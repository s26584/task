�csklearn.ensemble._forest
RandomForestClassifier
q )�q}q(X   base_estimatorqcsklearn.tree._classes
DecisionTreeClassifier
q)�q}q(X	   criterionqX   giniqX   splitterq	X   bestq
X	   max_depthqNX   min_samples_splitqKX   min_samples_leafqKX   min_weight_fraction_leafqG        X   max_featuresqNX   max_leaf_nodesqNX   random_stateqNX   min_impurity_decreaseqG        X   class_weightqNX	   ccp_alphaqG        X   _sklearn_versionqX   1.0.2qubX   n_estimatorsqKX   estimator_paramsq(hhhhhhhhhhtqX	   bootstrapq�X	   oob_scoreq�X   n_jobsqNhK X   verboseqK X
   warm_startq�hNX   max_samplesqNhhhNhKhKhG        hX   autoq hNhG        hG        X   feature_names_in_q!cnumpy.core.multiarray
_reconstruct
q"cnumpy
ndarray
q#K �q$Cbq%�q&Rq'(KK�q(cnumpy
dtype
q)X   O8q*���q+Rq,(KX   |q-NNNJ����J����K?tq.b�]q/(X   Ageq0X	   RestingBPq1X   Cholesterolq2X	   FastingBSq3X   MaxHRq4X   Oldpeakq5X   Mq6X   ATAq7X   NAPq8X   TAq9X   Normalq:X   STq;X   Yq<X   Flatq=X   Upq>etq?bX   n_features_in_q@KX
   n_outputs_qAKX   classes_qBh"h#K �qCh%�qDRqE(KK�qFh)X   i8qG���qHRqI(KX   <qJNNNJ����J����K tqKb�C               qLtqMbX
   n_classes_qNKX   base_estimator_qOhX   estimators_qP]qQ(h)�qR}qS(hhh	h
hNhKhKhG        hh hNhJ�
hG        hNhG        h@KhAKhBh"h#K �qTh%�qURqV(KK�qWh)X   f8qX���qYRqZ(KhJNNNJ����J����K tq[b�C              �?q\tq]bhNcnumpy.core.multiarray
scalar
q^hIC       q_�q`RqaX   max_features_qbKX   tree_qccsklearn.tree._tree
Tree
qdKh"h#K �qeh%�qfRqg(KK�qhhI�C       qitqjbK�qkRql}qm(hKX
   node_countqnK�X   nodesqoh"h#K �qph%�qqRqr(KKυqsh)X   V56qt���quRqv(Kh-N(X
   left_childqwX   right_childqxX   featureqyX	   thresholdqzX   impurityq{X   n_node_samplesq|X   weighted_n_node_samplesq}tq~}q(hwh)X   i8q����q�Rq�(KhJNNNJ����J����K tq�bK �q�hxh�K�q�hyh�K�q�hzhZK�q�h{hZK �q�h|h�K(�q�h}hZK0�q�uK8KKtq�b�BH-         t                    �?h�|�`�?�           ��@                          Pe@(4w%��?�            �w@                           �? ��+,��?O            @_@                           W@p��%���?+            @Q@                           �?      �?              @������������������������       �                     �?������������������������       �                     �?                           �?�����?)            �P@	       
       
             �?�i�y�?&            �O@������������������������       �        
             ,@                          @^@@9G��?            �H@                           �J@�r����?             .@������������������������       �                      @                           [@����X�?             @                          �W@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     A@                          �`@      �?             @                        `ff�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �        $             L@       i       	             �?B��T��?�            p@       Z                    �?�\����?�            �n@       5                    �?|g�&��?�            `i@       (                   @q@�\��N��?             C@       #                    a@�q�q�?	             (@                            b@      �?              @������������������������       �                     @!       "                    �?      �?             @������������������������       �                     �?������������������������       �                     @$       '                    �?      �?             @%       &                    @J@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @)       4                    �?�n_Y�K�?             :@*       3                   �b@�G��l��?             5@+       0                   @e@d}h���?	             ,@,       /                    @I@ףp=
�?             $@-       .                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @1       2                   u@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     @6       W                    �?d#,����?k            �d@7       V                    �?�O��e�?b            �b@8       9                    �?�t`�4 �?O            �^@������������������������       �                     0@:       C                    �F@����&��?D            �Z@;       B                   Xp@X�Cc�?	             ,@<       A                    @X�<ݚ�?             "@=       >                     C@z�G�z�?             @������������������������       �                      @?       @                    _@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @D       U                    �L@���.�6�?;             W@E       P                    @L@\#r��?%            �N@F       O                    �?`'�J�?             �I@G       H       
             �?�nkK�?             G@������������������������       �                      @I       J                    `@���7�?             F@������������������������       �                     >@K       L                   �p@؇���X�?             ,@������������������������       �                     &@M       N                   Pt@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @Q       R       
             �?���Q��?             $@������������������������       �                     @S       T                   @[@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     ?@������������������������       �                     <@X       Y                    m@z�G�z�?	             .@������������������������       �                     @������������������������       �                     (@[       \                     F@����X�?             E@������������������������       �                      @]       h                   @q@�t����?             A@^       _                   �[@�C��2(�?            �@@������������������������       �                     �?`       a                    �?      �?             @@������������������������       �                     �?b       c                    n@�g�y��?             ?@������������������������       �                     5@d       g                 ����?ףp=
�?             $@e       f                   0c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?j       k                    �?      �?
             (@������������������������       �                     @l       m                   0l@�q�q�?             "@������������������������       �                      @n       s                    �?؇���X�?             @o       r                    �?�q�q�?             @p       q                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @u       �                    �?��p
,�?�             s@v       �                    �?�gc� �?�             o@w       �                    @Lő����?�            `j@x       �                 pff�?X��J��?�             j@y       �                   �b@P���Q�?q            �f@z       �                    @N@ �Jj�G�?h            �d@{       �       
             �? YyH9�?`            �b@|       }                    �?��<b�ƥ?             G@������������������������       �                     4@~       �                    �? ��WV�?             :@       �                   �\@@4և���?	             ,@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@������������������������       �                     (@������������������������       �        E            @Z@�       �                 ����?؇���X�?             ,@�       �                    �?����X�?             @�       �                   �_@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �       
             �?���Q��?	             .@�       �                    �?և���X�?             @������������������������       �                      @�       �                   �m@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    �?      �?              @������������������������       �                     @�       �                    �?���Q��?             @�       �                   @k@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                    �?V�a�� �?             =@�       �                    �?���!pc�?             6@������������������������       �                     &@�       �                   p`@�eP*L��?             &@������������������������       �                     @�       �                   @k@����X�?             @�       �                   �b@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                      @�       �                   �X@P����?             C@������������������������       �                      @�       �                    �?<ݚ)�?             B@�       �                   0a@r�q��?             >@�       �                     L@�t����?             1@������������������������       �                     $@�       �                   �`@����X�?             @�       �                 ����?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                     N@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     *@������������������������       �                     @�       �                    �?���b���?             �L@�       �                    �?�q�q�?             H@�       �                    �?��Hg���?            �F@�       �                    �?<ݚ)�?             B@�       �                   Pd@�û��|�?             7@�       �                   �_@     ��?
             0@�       �                     P@      �?             @������������������������       �                      @������������������������       �                      @�       �                   �b@�8��8��?             (@������������������������       �                      @�       �                   �p@      �?             @������������������������       �                     @������������������������       �                     �?�       �                   Pe@؇���X�?             @������������������������       �                     @�       �                   pf@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   @a@8�Z$���?             *@������������������������       �                     $@�       �       
             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     "@������������������������       �                     @������������������������       �                     "@q�tq�bX   valuesq�h"h#K �q�h%�q�Rq�(KK�KK�q�hZ�B�       �r@     �x@      K@     �t@      @     @^@      @     @P@      �?      �?              �?      �?              @      P@       @     �N@              ,@       @     �G@       @      *@               @       @      @       @       @               @       @                      @              A@      �?      @      �?      �?              �?      �?                       @              L@      I@     �i@      F@      i@      @@     `e@      2@      4@       @      @      @      �?      @              @      �?              �?      @              �?      @      �?      �?      �?                      �?               @      $@      0@      $@      &@      @      &@      �?      "@      �?      �?              �?      �?                       @       @       @               @       @              @                      @      ,@     �b@      &@     `a@      &@     �[@              0@      &@     �W@      @      "@      @      @      �?      @               @      �?       @               @      �?              @                      @      @     �U@      @     �K@       @     �H@       @      F@               @       @      E@              >@       @      (@              &@       @      �?       @                      �?              @      @      @              @      @       @               @      @                      ?@              <@      @      (@      @                      (@      (@      >@       @              @      >@      @      >@      �?               @      >@      �?              �?      >@              5@      �?      "@      �?      �?      �?                      �?               @      �?              @      @      @              @      @       @              �?      @      �?       @      �?      �?              �?      �?                      �?              @     @n@      P@     `k@      >@     @h@      1@     @h@      .@     `e@      "@     @d@      @     �b@      �?     �F@      �?      4@              9@      �?      *@      �?      �?      �?              �?      �?              (@              (@             @Z@              (@       @      @       @      �?       @      �?                       @      @              @              "@      @      @      @       @              �?      @              @      �?              @       @      @              @       @      �?       @      �?                       @       @              7@      @      0@      @      &@              @      @              @      @       @      �?       @      �?                       @      @              @                       @      9@      *@               @      9@      &@      9@      @      (@      @      $@               @      @      �?      �?      �?                      �?      �?      @              @      �?              *@                      @      7@      A@      ,@      A@      &@      A@      &@      9@      "@      ,@      @      *@       @       @       @                       @      �?      &@               @      �?      @              @      �?              @      �?      @              �?      �?              �?      �?               @      &@              $@       @      �?              �?       @                      "@      @              "@        q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJ/��hG        hNhG        h@KhAKhBh"h#K �q�h%�q�Rq�(KK�q�hZ�C              �?q�tq�bhNh^hIC       q��q�Rq�hbKhchdKh"h#K �q�h%�q�Rq�(KK�q�hI�C       q�tq�bK�q�Rq�}q�(hKhnK�hoh"h#K �q�h%�q�Rq�(KKǅq�hv�B�+         ~                    �?�ٳU=��?�           ��@       =                    �?R���Q�?�             y@       (                   �c@�&z{�?^            �c@                          �a@Riv����?H             ]@                           �L@����?�?            �F@                           �?���7�?             6@������������������������       �                     3@       	                    ��q�q�?             @������������������������       �                     �?
                          �Z@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     7@                           �?v���EO�?.            �Q@                          �^@�G�z��?             4@������������������������       �                      @                           `P@      �?             (@                          �`@ףp=
�?             $@                        ����?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                      @       !                 ����?�t����?"            �I@                          �k@д>��C�?             =@                           �?      �?              @������������������������       �                     @������������������������       �                     @                          �p@���N8�?             5@������������������������       �                     *@                            �?      �?              @������������������������       �                     �?������������������������       �                     @"       #                    �N@���7�?             6@������������������������       �        
             ,@$       %                   `a@      �?              @������������������������       �                     @&       '       
             �?      �?             @������������������������       �                     @������������������������       �                     �?)       .                    �?�p ��?            �D@*       +                   �`@�r����?             .@������������������������       �                     (@,       -                   �`@�q�q�?             @������������������������       �                      @������������������������       �                     �?/       4                    @I@R�}e�.�?             :@0       3                    �?��S�ۿ?             .@1       2                    @E@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     (@5       6                    �?�eP*L��?             &@������������������������       �                      @7       8                    ]@�q�q�?             "@������������������������       �                      @9       <                    �?؇���X�?             @:       ;                    X@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @>       }                    �R@,�!�?�            `n@?       j                    �L@�l�T{�?�             n@@       A                   �U@��ϻ�r�?W            ``@������������������������       �                      @B       e                   �e@�����?V             `@C       N                    �?����y7�?S            @_@D       I                   �l@������?             1@E       H                   `a@      �?             @F       G                     I@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @J       M                    ]@$�q-�?             *@K       L                   �Z@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     "@O       d                 ����?�>����?G             [@P       a                    �?      �?*             P@Q       `                   �l@lGts��?#            �K@R       S       
             �?b�h�d.�?            �A@������������������������       �                     "@T       Y                    �?�θ�?             :@U       V                    �J@�KM�]�?             3@������������������������       �        	             0@W       X                    �K@�q�q�?             @������������������������       �                      @������������������������       �                     �?Z       [                   �`@և���X�?             @������������������������       �                      @\       _                   �_@z�G�z�?             @]       ^                   �j@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     4@b       c                    �G@�<ݚ�?             "@������������������������       �                      @������������������������       �                     @������������������������       �                     F@f       i                   �g@      �?             @g       h                   u@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?k       l                    �?h㱪��?I            �[@������������������������       �        
             1@m       n                   �j@H��2�??            @W@������������������������       �                    �C@o       p                    @N@�>����?%             K@������������������������       �        	             ,@q       r                    �?ףp=
�?             D@������������������������       �                     @s       z                    �?(N:!���?            �A@t       y                   �Z@(;L]n�?             >@u       x                   `a@؇���X�?             @v       w       
             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     7@{       |                    �P@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @       �                    �K@F��ӭ��?�             r@�       �                 ����?���\��?z            �h@�       �                    �?x�@�E-�?f             d@�       �                   �h@��K˱F�?]            �a@�       �                    �?�KM�]�?             C@�       �                    @F@؇���X�?             <@�       �                    �?�q�q�?             (@�       �                    ]@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     0@������������������������       �                     $@�       �       
             �?@��!�Q�?D            @Z@������������������������       �                     A@�       �                    @D@ ��PUp�?0            �Q@�       �                   �f@$�q-�?
             *@������������������������       �        	             (@������������������������       �                     �?������������������������       �        &             M@�       �                    `@r�q��?	             2@������������������������       �                     @������������������������       �                     .@�       �                    d@�\��N��?             C@������������������������       �                     @�       �                   `b@f���M�?             ?@�       �                    �?r�q��?             8@�       �                   �_@      �?             (@�       �                   c@և���X�?             @������������������������       �                      @�       �                    �E@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                   �`@�q�q�?             (@������������������������       �                     @�       �                   pi@�����H�?             "@������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                   �O@���R��?8            @V@�       �                    �?"pc�
�?             6@�       �                    �?������?             .@�       �                   �`@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     $@������������������������       �                     @�       �                    �?�#}7��?+            �P@�       �                    �?�C��2(�?             6@�       �                    �N@���N8�?             5@�       �                    `@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �        
             1@������������������������       �                     �?�       �                    �?��S���?            �F@�       �                   �`@���B���?             :@�       �                   ``@�eP*L��?             &@�       �                   �a@      �?              @������������������������       �                     @�       �                   �^@      �?             @������������������������       �                     �?�       �                   �_@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     .@�       �                   �d@�S����?
             3@�       �                    �L@�����H�?	             2@������������������������       �                      @������������������������       �                     0@������������������������       �                     �?q�tq�bh�h"h#K �q�h%�q�Rq�(KK�KK�q�hZ�Bp       �q@     py@      N@     @u@      C@     �]@      2@     �X@      �?      F@      �?      5@              3@      �?       @              �?      �?      �?      �?                      �?              7@      1@      K@      &@      "@       @              @      "@      �?      "@      �?      @              @      �?                      @       @              @     �F@      @      8@      @      @              @      @              �?      4@              *@      �?      @      �?                      @      �?      5@              ,@      �?      @              @      �?      @              @      �?              4@      5@      *@       @      (@              �?       @               @      �?              @      3@      �?      ,@      �?       @      �?                       @              (@      @      @               @      @      @               @      @      �?      @      �?              �?      @              @              6@     �k@      4@     �k@      0@     �\@       @              ,@     �\@      (@     @\@      @      *@      @      �?      �?      �?              �?      �?               @              �?      (@      �?      @              @      �?                      "@       @      Y@       @      L@      @     �H@      @      =@              "@      @      4@       @      1@              0@       @      �?       @                      �?      @      @               @      @      �?       @      �?       @                      �?       @                      4@       @      @       @                      @              F@       @       @       @      �?              �?       @                      �?      @     �Z@              1@      @     @V@             �C@      @      I@              ,@      @      B@              @      @      ?@      �?      =@      �?      @      �?       @               @      �?                      @              7@      @       @      @                       @       @             �k@     �P@     �e@      :@      c@       @     @a@      @      A@      @      8@      @       @      @      �?      @              @      �?              @              0@              $@              Z@      �?      A@             �Q@      �?      (@      �?      (@                      �?      M@              .@      @              @      .@              4@      2@              @      4@      &@      *@      &@      "@      @      @      @       @               @      @       @                      @      @              @       @      @              �?       @      �?                       @      @              H@     �D@      @      2@      @      &@      @      �?              �?      @                      $@              @      F@      7@      4@       @      4@      �?      @      �?      @                      �?      1@                      �?      8@      5@      5@      @      @      @      @       @      @               @       @      �?              �?       @               @      �?                      @      .@              @      0@       @      0@       @                      0@      �?        q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJu�7hG        hNhG        h@KhAKhBh"h#K �q�h%�q�Rq�(KK�q�hZ�C              �?q�tq�bhNh^hIC       q��q�Rq�hbKhchdKh"h#K �q�h%�q�Rq�(KK�q�hI�C       q�tq�bK�q�Rq�}q�(hKhnK�hoh"h#K �q�h%�q�Rq�(KKՅq�hv�B�.         `                    �?�����?�           ��@       K                    �?t�I��n�?�            �u@       >                    �?��e2A�?�             q@       %                    �?r�qG�?|             h@              
             �? ���g=�?Z            @a@       	                    �?z�G�z�?$            �K@                          e@���N8�?             5@������������������������       �                     �?������������������������       �                     4@
                          �q@�t����?             A@                          Pf@d}h���?             <@                        ����?և���X�?             @                          pc@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @                           @�����?             5@������������������������       �                     3@������������������������       �                      @                           a@�q�q�?             @������������������������       �                     �?                          �_@z�G�z�?             @������������������������       �                     @������������������������       �                     �?       $                   �b@ ,U,?��?6            �T@                        833�?�[|x��?+            �O@                          d@ 7���B�?$             K@������������������������       �                     @@                          @d@�C��2(�?             6@������������������������       �                      @������������������������       �                     4@        !                    @F@�q�q�?             "@������������������������       �                     @"       #                 ����?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     4@&       9                   n@�q�q�?"             K@'       0                   `a@�D����?             E@(       -       
             �?8�Z$���?             :@)       *                    �?      �?              @������������������������       �                     @+       ,                   �a@���Q��?             @������������������������       �                     @������������������������       �                      @.       /                   @^@�����H�?
             2@������������������������       �                      @������������������������       �                     0@1       2                    �?     ��?	             0@������������������������       �                     @3       8                    �?�θ�?             *@4       5                    a@�C��2(�?             &@������������������������       �                     @6       7                 033�?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @:       =                    a@�8��8��?	             (@;       <                    �L@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @?       F                 ����?��Y��]�?;            �T@@       A                    c@�k~X��?3             R@������������������������       �        /             Q@B       C                    �K@      �?             @������������������������       �                      @D       E                   `c@      �?              @������������������������       �                     �?������������������������       �                     �?G       J                 pff�?ףp=
�?             $@H       I                   p`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @L       Q                    �?�eP*L��?,            @S@M       N                    �F@      �?             0@������������������������       �                     �?O       P                   �r@��S�ۿ?
             .@������������������������       �        	             ,@������������������������       �                     �?R       S                   �O@N1���?!            �N@������������������������       �        
             5@T       _       
             �?z�G�z�?             D@U       ^                    �?�X����?             6@V       ]                 ����?�q�q�?             (@W       X                   0b@r�q��?             @������������������������       �                     @Y       Z                    �?�q�q�?             @������������������������       �                     �?[       \                   �`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     $@������������������������       �                     2@a       �                   �a@<ܹ���?�            u@b       m                   `h@���m��?�            �n@c       l                    �?��Y��]�?4            �T@d       k                   @_@��S�ۿ?             >@e       f                   �]@z�G�z�?             $@������������������������       �                     @g       j                    �?���Q��?             @h       i                    X@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �        	             4@������������������������       �        $             J@n       �                    �?���Ȓ��?h            `d@o       v                   `[@�*/�8V�?V            �a@p       u                 433�?����?�?            �F@q       r                   0o@@4և���?             ,@������������������������       �                     (@s       t                   �Y@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     ?@w       �                    �?8��8���?=             X@x       y                    �D@և���X�?             ,@������������������������       �                     @z       �                    �?���Q��?             $@{       ~                    �?X�<ݚ�?             "@|       }                     P@�q�q�?             @������������������������       �                      @������������������������       �                     �?       �                    �J@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     �?�       �                    �J@������?5            �T@�       �                   `j@H�V�e��?             A@�       �                   pa@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �?�חF�P�?             ?@�       �                    �?HP�s��?             9@�       �                   hq@r�q��?             (@������������������������       �                     @�       �                   ``@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �        	             *@�       �                     H@      �?             @������������������������       �                     �?�       �                    @���Q��?             @�       �                   �`@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                 ����?@��8��?             H@�       �                    �L@�X�<ݺ?             2@�       �                   `_@؇���X�?             @������������������������       �                     @�       �                   Pq@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@������������������������       �                     >@�       �                    @M@�GN�z�?             6@������������������������       �                      @�       �                   �j@X�Cc�?             ,@������������������������       �                     @�       �                 ����?"pc�
�?             &@�       �                    �P@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                    �?�y�ʍ+�??             W@�       �                    �?���N8�?             5@�       �       	             �?��S�ۿ?             .@������������������������       �                     ,@������������������������       �                     �?�       �                    �?�q�q�?             @�       �                    �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?�       �                    �?���BK�?2            �Q@�       �                     O@�&!��?            �E@�       �                    �M@��Q��?             D@�       �                   �?j���� �?             A@������������������������       �                     $@�       �                    �I@�q�q�?             8@�       �                   �d@�q�q�?
             (@�       �                   �a@      �?              @������������������������       �                     �?������������������������       �                     @�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @�       �                   �p@r�q��?             (@�       �                    m@ףp=
�?             $@�       �                   `d@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                   0r@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �?@4և���?             <@�       �                     M@ ��WV�?             :@������������������������       �                     4@�       �                   �_@r�q��?             @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �n@      �?              @������������������������       �                     �?������������������������       �                     �?q�tq�bh�h"h#K �q�h%�q�Rq�(KK�KK�q�hZ�BP       �s@     �w@     �o@      X@     �k@      K@     �a@      J@     �^@      0@      F@      &@      4@      �?              �?      4@              8@      $@      6@      @      @      @      @       @      @                       @               @      3@       @      3@                       @       @      @      �?              �?      @              @      �?             �S@      @      M@      @      J@       @      @@              4@       @               @      4@              @      @      @               @      @              @       @              4@              2@      B@      1@      9@      @      6@       @      @              @       @      @              @       @               @      0@       @                      0@      *@      @      @              $@      @      $@      �?      @              @      �?      @                      �?               @      �?      &@      �?      @      �?                      @               @      T@       @     �Q@      �?      Q@              @      �?       @              �?      �?              �?      �?              "@      �?      �?      �?              �?      �?               @             �A@      E@       @      ,@      �?              �?      ,@              ,@      �?             �@@      <@              5@     �@@      @      .@      @      @      @      @      �?      @               @      �?      �?              �?      �?      �?                      �?              @      $@              2@             �L@     �q@      6@     �k@       @      T@       @      <@       @       @              @       @      @       @      �?              �?       @                       @              4@              J@      4@     �a@      .@     �_@      �?      F@      �?      *@              (@      �?      �?              �?      �?                      ?@      ,@     �T@      @       @              @      @      @      @      @       @      �?       @                      �?      @      @      @                      @      �?               @     �R@      @      ;@       @      �?       @                      �?      @      :@       @      7@       @      $@              @       @      @              @       @                      *@      @      @      �?               @      @       @      �?       @                      �?               @      �?     �G@      �?      1@      �?      @              @      �?      �?      �?                      �?              &@              >@      @      1@               @      @      "@      @               @      "@       @       @       @                       @              @     �A@     �L@      0@      @      ,@      �?      ,@                      �?       @      @       @      @              @       @                      �?      3@      J@      1@      :@      ,@      :@      ,@      4@              $@      ,@      $@      @       @      �?      @      �?                      @      @      �?              �?      @              $@       @      "@      �?      @      �?      @                      �?      @              �?      �?              �?      �?                      @      @               @      :@      �?      9@              4@      �?      @              @      �?       @      �?                       @      �?      �?      �?                      �?q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJ��!XhG        hNhG        h@KhAKhBh"h#K �q�h%�q�Rq�(KK�q�hZ�C              �?q�tq�bhNh^hIC       q݆q�Rq�hbKhchdKh"h#K �q�h%�q�Rq�(KK�q�hI�C       q�tq�bK�q�Rq�}q�(hKhnK�hoh"h#K �q�h%�q�Rq�(KKӅq�hv�B(.         �                    �?�կZ���?�           ��@       y                    �?�� ƞ��?i           P�@       h                   �c@���T�(�?            y@       %                 033�?�	����?�            0v@                          �a@������?N            @]@                           �?�+��<��?;            �U@                        ����?��� ��?             ?@                           �? 	��p�?             =@	                          �e@ףp=
�?             4@
              
             �?�q�q�?             @������������������������       �                     �?                           P@z�G�z�?             @                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     ,@������������������������       �                     "@������������������������       �                      @                        833�?z�G�z�?$            �K@������������������������       �                    �C@                           �?     ��?
             0@                          �`@8�Z$���?             *@������������������������       �                     @                          `m@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @       $                    �?�חF�P�?             ?@                           �?��<b���?             7@������������������������       �                     @        !                    �?�}�+r��?             3@������������������������       �                     &@"       #                     K@      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                      @&       ?                    �?  6�W �?�            �m@'       4                 ����?`�Q��?%             I@(       -                   Pn@     ��?             0@)       ,                    �?r�q��?             @*       +                    �N@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @.       3       
             �?z�G�z�?             $@/       0                     K@���Q��?             @������������������������       �                      @1       2                    �L@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @5       >                    �?H�V�e��?             A@6       9                    �?p�ݯ��?             3@7       8                   `c@����X�?             @������������������������       �                     @������������������������       �                      @:       =                 ���@r�q��?
             (@;       <                    �?����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     .@@       A                   �U@��`ۻ��?x            �g@������������������������       �                     �?B       e                    �R@C���?w            `g@C       ^                    �L@���.�6�?u             g@D       Q                   0i@�ʠ����?B            �Z@E       F       
             �?d}h���?             E@������������������������       �        	             .@G       H                   `_@�q�q�?             ;@������������������������       �                     &@I       P                    �?     ��?             0@J       K                    �?"pc�
�?             &@������������������������       �                     @L       M                    �C@����X�?             @������������������������       �                     �?N       O                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @R       W                    @G@��ɉ�?*            @P@S       V                   @n@ףp=
�?             $@T       U                    ^@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @X       Y                 033@ �Jj�G�?"            �K@������������������������       �                    �G@Z       ]       
             �?      �?              @[       \                 `ff@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @_       `                 033�?�e���@�?3            @S@������������������������       �                    �E@a       d                    �?г�wY;�?             A@b       c                   �b@ �q�q�?             8@������������������������       �                     7@������������������������       �                     �?������������������������       �                     $@f       g                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @i       r                   m@���Q��?            �F@j       q                   �^@�X����?             6@k       p                    @L@�z�G��?             $@l       o                    �E@�<ݚ�?             "@m       n                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �        	             (@s       x                    �?�LQ�1	�?             7@t       u                    �?���N8�?             5@������������������������       �        	             3@v       w                 @33�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @z       �                    �?8�A�0��?b            @c@{       �       
             �?ȵHPS!�?6            �S@|                          `d@�θ�?             :@}       ~                 @33�?z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                   pe@�����?             5@������������������������       �                     0@�       �                    �?���Q��?             @������������������������       �                     �?�       �                   �l@      �?             @������������������������       �                      @������������������������       �                      @�       �                   �O@0G���ջ?$             J@�       �                 ����?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �G@�       �                   ``@p9W��S�?,             S@�       �                   �c@�s��:��?             C@�       �                    �?��H�}�?             9@�       �                    �Q@8�A�0��?             6@�       �                    �?�G�z��?             4@������������������������       �                      @�       �                   `]@b�2�tk�?             2@������������������������       �                     @�       �                    ����|���?             &@������������������������       �                     �?�       �                 ����?�z�G��?             $@������������������������       �                      @�       �                    �O@      �?              @�       �                   �l@����X�?             @�       �       
             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    ]@$�q-�?             *@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@�       �                 tff�?P�Lt�<�?             C@�       �                 ����?�8��8��?             (@������������������������       �                     &@������������������������       �                     �?������������������������       �                     :@�       �                   �^@t�U����?X            �`@�       �                    �?      �?             0@������������������������       �                     @�       �       
             �?z�G�z�?             $@�       �                   0a@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                    c@ ,��-�?M            �]@�       �                    �? '��h�?F            @[@�       �                    �?p�qG�?;             X@�       �                 ����?�J�4�?             9@������������������������       �                     $@�       �                   �\@������?             .@������������������������       �                      @�       �                   @b@8�Z$���?             *@������������������������       �                     @�       �       
             �?����X�?             @�       �                 ����?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �K@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    �? ��PUp�?/            �Q@������������������������       �                     6@�       �                   �a@@�E�x�?!            �H@�       �                 @33�?      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                    �D@������������������������       �                     *@�       �                    �?�q�q�?             "@������������������������       �                     �?�       �                    @K@      �?              @������������������������       �                     @�       �                   �b@      �?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @q�tq�bh�h"h#K �q�h%�q�Rq�(KK�KK�q�hZ�B0       `s@     �w@      h@     �v@     @Y@     �r@     �R@     �q@     �E@     �R@      C@      H@      ;@      @      ;@       @      2@       @      @       @              �?      @      �?       @      �?       @                      �?       @              ,@              "@                       @      &@      F@             �C@      &@      @      &@       @      @              @       @      @                       @              @      @      :@      @      2@      @              �?      2@              &@      �?      @      �?                      @               @      ?@     �i@      0@      A@      "@      @      �?      @      �?      �?              �?      �?                      @       @       @      @       @       @              �?       @               @      �?              @              @      ;@      @      (@      @       @      @                       @       @      $@       @      @              @       @                      @              .@      .@     �e@      �?              ,@     �e@      (@     �e@      &@      X@      "@     �@@              .@      "@      2@              &@      "@      @      "@       @      @              @       @              �?      @      �?      @                      �?              @       @     �O@      �?      "@      �?      �?      �?                      �?               @      �?      K@             �G@      �?      @      �?      @      �?                      @              @      �?      S@             �E@      �?     �@@      �?      7@              7@      �?                      $@       @      �?              �?       @              ;@      2@      @      .@      @      @      @       @       @       @               @       @              @                      �?              (@      4@      @      4@      �?      3@              �?      �?              �?      �?                       @     �V@     �O@     @Q@      "@      4@      @      �?      @      �?                      @      3@       @      0@              @       @      �?               @       @               @       @             �H@      @       @      @       @                      @     �G@              6@      K@      5@      1@      "@      0@      "@      *@      "@      &@       @              @      &@              @      @      @              �?      @      @       @              @      @      @       @      �?       @               @      �?              @                      �?               @              @      (@      �?      �?      �?      �?                      �?      &@              �?     �B@      �?      &@              &@      �?                      :@     �]@      0@       @       @              @       @       @       @       @       @                       @      @             �[@       @      Z@      @     �V@      @      5@      @      $@              &@      @               @      &@       @      @              @       @      �?      �?      �?                      �?      @      �?      @                      �?     �Q@      �?      6@              H@      �?      @      �?      @                      �?     �D@              *@              @      @      �?              @      @      @              �?      @      �?      �?      �?                      �?               @q�tq�bubhhubh)�q�}q�(hhh	h
hNhKhKhG        hh hNhJC�NhG        hNhG        h@KhAKhBh"h#K �q�h%�q�Rq�(KK�q�hZ�C              �?q�tq�bhNh^hIC       q��q�Rq�hbKhchdKh"h#K �r   h%�r  Rr  (KK�r  hI�C       r  tr  bK�r  Rr  }r  (hKhnK�hoh"h#K �r	  h%�r
  Rr  (KKۅr  hv�B�/         �                    �?�T�%y��?�           ��@       E                    �?`�'�?
           �x@                          `[@�&|�&��?�            �p@                           �?     ��?             0@������������������������       �                     @������������������������       �                     *@       ,                    @L@Ί�C�o�?�            �o@                          �`@(l58��?�            �h@	       
                   �\@��Hg���?            �F@������������������������       �                      @                           �?V������?            �B@                           �?� �	��?             9@              
             �?d}h���?             ,@������������������������       �                      @                           �?�8��8��?             (@������������������������       �                     &@������������������������       �                     �?������������������������       �        	             &@������������������������       �                     (@                          0c@�C��2(�?k            @c@������������������������       �        $             H@       !                    ]@^�!~X�?G            �Z@                          @[@�X����?             6@������������������������       �                     &@                            �?���|���?
             &@                           �?�<ݚ�?             "@                          �l@      �?              @������������������������       �                     @                          0f@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @"       #                    �?�8��8��?5             U@������������������������       �                     8@$       +                    �?�?�P�a�?'             N@%       &                   �j@��G���?            �B@������������������������       �                     1@'       *                   @b@��Q��?             4@(       )                   �d@�E��ӭ�?             2@������������������������       �                     @������������������������       �                     *@������������������������       �                      @������������������������       �                     7@-       8                    �?�q����?%            �J@.       /                   �c@���Q��?             .@������������������������       �                     @0       1                    �?�eP*L��?             &@������������������������       �                      @2       7                    �?X�<ݚ�?             "@3       6                    �?�q�q�?             @4       5                    b@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @9       :                   �O@>A�F<�?             C@������������������������       �                      @;       <                   �b@4?,R��?             B@������������������������       �                     7@=       D                    �?�n_Y�K�?	             *@>       ?                    �M@���!pc�?             &@������������������������       �                     @@       C                    �?���Q��?             @A       B       
             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                      @F       {                    �?4�.�A�?S            �_@G       p                    �?r�qG�?>             X@H       c                    �?^��4m�?-            �R@I       \                   0c@���*�?$             N@J       S                   �`@ȵHPS!�?             J@K       N                    �M@�>4և��?             <@L       M                 ����?����X�?	             ,@������������������������       �                     @������������������������       �                     $@O       P                   @_@@4և���?	             ,@������������������������       �                     "@Q       R                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @T       U                   �l@ �q�q�?             8@������������������������       �                     3@V       [       
             �?z�G�z�?             @W       X                   �a@�q�q�?             @������������������������       �                     �?Y       Z                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @]       ^                   �d@      �?              @������������������������       �                     @_       b                 ����?      �?             @`       a                   �e@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @d       k                   �^@և���X�?	             ,@e       f                   �\@r�q��?             @������������������������       �                     �?g       h       
             �?z�G�z�?             @������������������������       �                     @i       j                   �p@      �?              @������������������������       �                     �?������������������������       �                     �?l       m                    @L@      �?              @������������������������       �                     @n       o                   �^@      �?              @������������������������       �                     �?������������������������       �                     �?q       v                    �?�X����?             6@r       u                    a@�<ݚ�?             2@s       t                   �^@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �        	             (@w       z                    �?      �?             @x       y                    ]@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?|       �                   �c@���Q��?             >@}       �                    �?j���� �?             1@~       �                    �?      �?             0@       �                 `ff�?��
ц��?
             *@�       �                   ph@      �?              @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     �?�       �                    �L@8�Z$���?	             *@������������������������       �                     &@������������������������       �                      @�       �                   �h@8�ǫ�0�?�            `r@�       �                    �? ѯ��?D            �Z@�       �                   �_@�8��8��?.             R@������������������������       �                     G@�       �                   �U@�θ�?             :@������������������������       �                     �?�       �                    �?z�G�z�?             9@�       �                    @G@�S����?             3@�       �                    `@      �?              @������������������������       �                      @�       �       
             �?r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     &@�       �                    �?�q�q�?             @�       �                    �?�q�q�?             @�       �                   Pa@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                    �A@�       �                   �b@p�~;��?y            `g@�       �                    �?�S�%3��?k            �c@�       �                   �[@������?b             b@�       �                    �K@և���X�?             @�       �                    @G@�q�q�?             @�       �       
             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �       
             �?D��*�4�?]            @a@�       �                    �L@      �?)             P@�       �                    @L@�>����?             ;@�       �                   �\@�nkK�?             7@�       �                   �[@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     4@�       �                 033�?      �?             @�       �                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                    �B@�       �                 ����?������?4            �R@�       �                    �? �o_��?             9@�       �                   @m@�����H�?             "@������������������������       �                     �?������������������������       �                      @�       �                   �k@      �?             0@������������������������       �                      @�       �                    @K@և���X�?             ,@������������������������       �                     @�       �                   `c@      �?              @������������������������       �                     @������������������������       �                      @�       �                    �?@�E�x�?#            �H@�       �                   �c@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                    �D@�       �                    �?X�Cc�?	             ,@�       �                   �_@�eP*L��?             &@������������������������       �                     @�       �                   `a@����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                   Pe@��X��?             <@�       �                   �i@      �?             8@������������������������       �                     "@�       �                    a@���Q��?	             .@������������������������       �                     @�       �                    �?�eP*L��?             &@������������������������       �                     @�       �                   0p@      �?              @������������������������       �                     @������������������������       �                      @�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @r  tr  bh�h"h#K �r  h%�r  Rr  (KK�KK�r  hZ�B�       �s@     pw@     �p@      `@     �j@      K@      @      *@      @                      *@     `j@     �D@     �e@      9@      A@      &@       @              :@      &@      ,@      &@      @      &@       @              �?      &@              &@      �?              &@              (@             �a@      ,@      H@              W@      ,@      .@      @      &@              @      @       @      @      �?      @              @      �?      �?              �?      �?              �?               @             @S@      @      8@             �J@      @      >@      @      1@              *@      @      *@      @              @      *@                       @      7@             �B@      0@      @      "@              @      @      @       @              @      @      @       @      @      �?      @                      �?              �?              @      ?@      @               @      ?@      @      7@               @      @       @      @      @               @      @       @      �?              �?       @                       @               @      J@     �R@      A@      O@      3@     �K@      &@     �H@      @      G@      @      7@      @      $@      @                      $@      �?      *@              "@      �?      @      �?                      @      �?      7@              3@      �?      @      �?       @              �?      �?      �?      �?                      �?               @      @      @      @              �?      @      �?      �?              �?      �?                       @       @      @      �?      @              �?      �?      @              @      �?      �?              �?      �?              @      �?      @              �?      �?              �?      �?              .@      @      ,@      @       @      @       @                      @      (@              �?      @      �?       @      �?                       @              �?      2@      (@      @      $@      @      $@      @      @      @       @               @      @                      @              @      �?              &@       @      &@                       @     �G@     �n@      @     @Y@      @     �P@              G@      @      4@      �?              @      4@      @      0@      @      @       @              �?      @      �?                      @              &@       @      @       @      �?      �?      �?      �?                      �?      �?                      @             �A@     �D@     @b@      6@      a@      *@     �`@      @      @       @      @       @      �?       @                      �?              @      �?              $@      `@       @      O@       @      9@      �?      6@      �?       @               @      �?                      4@      �?      @      �?      �?      �?                      �?               @             �B@       @     �P@      @      2@      �?       @      �?                       @      @      $@               @      @       @              @      @       @      @                       @      �?      H@      �?      @              @      �?                     �D@      "@      @      @      @      @               @      @              @       @              @              3@      "@      2@      @      "@              "@      @      @              @      @      @               @      @              @       @              �?      @      �?                      @r  tr  bubhhubh)�r  }r  (hhh	h
hNhKhKhG        hh hNhJ�R�[hG        hNhG        h@KhAKhBh"h#K �r  h%�r  Rr  (KK�r  hZ�C              �?r  tr  bhNh^hIC       r  �r  Rr  hbKhchdKh"h#K �r   h%�r!  Rr"  (KK�r#  hI�C       r$  tr%  bK�r&  Rr'  }r(  (hKhnK�hoh"h#K �r)  h%�r*  Rr+  (KKۅr,  hv�B�/         �                    �?�hu0���?�           ��@       [                   �b@v���a�?�            �v@                          �b@\#r��?�            s@                           �?�Ń��̧?2             U@       
                   `X@@4և���?             <@       	                    �?z�G�z�?             $@                           �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     2@������������������������       �                      L@       ,                    �?x��6S�?�            �k@       %                    �?�*/�8V�?"            �G@       "       	             �?��G���?            �B@       !                   �a@��hJ,�?             A@                           (s@�q�q�?             8@                          �r@�t����?             1@                           �?      �?             0@                           �L@������?             .@                           `@���Q��?             $@                          @^@؇���X�?             @                           �?      �?             @������������������������       �                      @              
             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     $@#       $                   �q@�q�q�?             @������������������������       �                     �?������������������������       �                      @&       '       
             �?      �?             $@������������������������       �                     @(       )                    �?r�q��?             @������������������������       �                     @*       +                   �m@�q�q�?             @������������������������       �                      @������������������������       �                     �?-       >       
             �?���(`�?n            �e@.       /                    �?xdQ�m��?3            @T@������������������������       �                      @0       7                   �j@���;QU�?.            @R@1       6                    �?���y4F�?             3@2       3                   pi@      �?	             0@������������������������       �                     $@4       5                   �`@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @8       =                    _@@3����?#             K@9       :                    @J@�C��2(�?             &@������������������������       �                     @;       <                    �J@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                    �E@?       H                    �?d۬����?;            @W@@       G                    �?�q�q�?
             (@A       B                   @[@���|���?	             &@������������������������       �                     @C       D                 433�?      �?              @������������������������       �                      @E       F                   �a@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?I       Z                    �?�>����?1            @T@J       K                   �_@��(\���?0             T@������������������������       �                     ;@L       U                    �?���C��?             �J@M       P                 433�?�����?             E@N       O                    Y@      �?             @������������������������       �                     �?������������������������       �                     @Q       T                 ����?P�Lt�<�?             C@R       S                     F@�8��8��?	             (@������������������������       �                     �?������������������������       �                     &@������������������������       �                     :@V       Y                   �\@"pc�
�?             &@W       X                    �Q@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     �?\       a                    V@�q�q�?(             N@]       ^                   �_@ףp=
�?             $@������������������������       �                     @_       `                    @      �?             @������������������������       �                     @������������������������       �                     �?b       k                   �l@�q�����?              I@c       f                    �?������?
             .@d       e                    �?      �?              @������������������������       �                     �?������������������������       �                     �?g       h                   0g@�θ�?             *@������������������������       �                      @i       j                    �?�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?l       q                    �?<=�,S��?            �A@m       n       
             �?      �?             @������������������������       �                      @o       p                    �?      �?              @������������������������       �                     �?������������������������       �                     �?r       w                    �?�4�����?             ?@s       v                    �?�<ݚ�?             "@t       u                   Pp@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @x       �       	             �?��2(&�?             6@y       z                   �b@r�q��?
             2@������������������������       �                     �?{       �                    @C@�t����?	             1@|       }                   �o@�q�q�?             @������������������������       �                     �?~                            @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     ,@������������������������       �                     @�       �                    I@41L�>V�?�            0t@�       �                    �?���N8�?             E@�       �                   0f@HP�s��?             9@�       �                    �? �q�q�?             8@�       �                   �Y@r�q��?             @������������������������       �                     @�       �                   �^@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     2@������������������������       �                     �?�       �                 ����?��.k���?	             1@�       �                    �?�z�G��?             $@�       �                    @D@      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                    @؇���X�?             @�       �                     M@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �L@�n3�F��?�            �q@�       �       
             �?h�qVhԳ?�            �k@�       �                    �?����1�?+            @R@������������������������       �                     <@�       �                     I@���V��?            �F@�       �                   0f@��+7��?             7@�       �                    �?��
ц��?	             *@�       �                    �?      �?              @�       �       	             �?؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     $@�       �                    @K@���7�?             6@������������������������       �                     0@�       �                   b@r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                   �o@�}��L�?\            �b@������������������������       �        B            @[@�       �                    �?������?            �D@�       �                     I@      �?             @@������������������������       �                     4@�       �                    �J@r�q��?             (@������������������������       �                      @������������������������       �                     $@������������������������       �                     "@�       �       	             �?>n�T��?%             M@�       �                 833�?��WV��?!             J@�       �                    d@d}h���?             <@�       �       
             �?�����?             5@�       �                    �?      �?              @�       �                    �Q@�q�q�?             @�       �                    �?���Q��?             @�       �                   @a@�q�q�?             @�       �                   @n@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                   �^@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     *@�       �                 ����?և���X�?             @�       �                    �?�q�q�?             @�       �                   �_@�q�q�?             @������������������������       �                     �?�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                   pb@�q�q�?             8@�       �                   �c@��S�ۿ?	             .@������������������������       �                     *@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?�q�q�?             "@������������������������       �                     �?�       �                    @M@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     @r-  tr.  bh�h"h#K �r/  h%�r0  Rr1  (KK�KK�r2  hZ�B�       �s@     `w@     �K@     `s@      >@     0q@       @     �T@       @      :@       @       @       @      @              @       @                      @              2@              L@      <@      h@      (@     �A@      @      >@      @      =@      @      3@      @      (@      @      (@      @      &@      @      @      �?      @      �?      @               @      �?      �?      �?                      �?              @      @                      @              �?      �?                      @              $@       @      �?              �?       @              @      @              @      @      �?      @               @      �?       @                      �?      0@     �c@      @      S@               @      @      Q@      @      .@      @      (@              $@      @       @      @                       @              @      �?     �J@      �?      $@              @      �?      @      �?                      @             �E@      &@     �T@      @      @      @      @              @      @      @               @      @       @      @                       @      �?              @     �R@      @     �R@              ;@      @     �G@      @      C@      @      �?              �?      @              �?     �B@      �?      &@      �?                      &@              :@       @      "@       @      @              @       @                      @              �?      9@     �A@      �?      "@              @      �?      @              @      �?              8@      :@      &@      @      �?      �?      �?                      �?      $@      @               @      $@      �?      $@                      �?      *@      6@      @      �?       @              �?      �?              �?      �?              $@      5@      @       @       @       @               @       @              @              @      3@      @      .@      �?               @      .@       @      �?      �?              �?      �?      �?                      �?              ,@              @     0p@      P@      $@      @@       @      7@      �?      7@      �?      @              @      �?       @               @      �?                      2@      �?               @      "@      @      @      @      �?              �?      @                       @      �?      @      �?       @               @      �?                      @      o@      @@     �j@      "@     �P@      @      <@              C@      @      1@      @      @      @       @      @      �?      @              @      �?              �?              @              $@              5@      �?      0@              @      �?      @                      �?     �b@       @     @[@             �C@       @      >@       @      4@              $@       @               @      $@              "@             �A@      7@      =@      7@      6@      @      3@       @      @       @      @       @      @       @       @      �?      �?      �?      �?                      �?      �?              �?      �?      �?                      �?      �?               @              *@              @      @       @      @       @      �?      �?              �?      �?              �?      �?                      @      �?              @      1@      �?      ,@              *@      �?      �?      �?                      �?      @      @      �?              @      @              @      @              @        r3  tr4  bubhhubh)�r5  }r6  (hhh	h
hNhKhKhG        hh hNhJ�v}hG        hNhG        h@KhAKhBh"h#K �r7  h%�r8  Rr9  (KK�r:  hZ�C              �?r;  tr<  bhNh^hIC       r=  �r>  Rr?  hbKhchdKh"h#K �r@  h%�rA  RrB  (KK�rC  hI�C       rD  trE  bK�rF  RrG  }rH  (hKhnK�hoh"h#K �rI  h%�rJ  RrK  (KKӅrL  hv�B(.         �                    �?��1j	��?�           ��@       A                 033�?�"�&z�?X           8�@       &                    �?�!g��?�            �n@                           �?r�q��?R            @a@                          �X@@4և���?D             \@������������������������       �                      @                        pff�?�1�`jg�?C            �[@                          Xt@��s�n�?@             Z@	       
                    �?`�E���?<            @X@������������������������       �                     :@                           b@�J�T�?+            �Q@������������������������       �        $            �J@                        @33�?�����H�?             2@                          d@؇���X�?             ,@������������������������       �                     (@������������������������       �                      @������������������������       �                     @                        @33�?և���X�?             @                           @J@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     �?                          a@r�q��?             @������������������������       �                     �?������������������������       �                     @                           �?
j*D>�?             :@������������������������       �                     @                           h@
;&����?             7@������������������������       �                      @       %                    �O@������?	             .@       $                    b@8�Z$���?             *@        !                   �_@�8��8��?             (@������������������������       �                     @"       #                   �d@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                      @'       6                   �b@�iʫ{�?A            �Z@(       -                    �?����"$�?3            �U@)       *                   �`@�q�q�?             "@������������������������       �                     @+       ,                   �?���Q��?             @������������������������       �                     @������������������������       �                      @.       5                    �?�e���@�?,            @S@/       0                   @l@����?�?            �F@������������������������       �                     ?@1       4                    \@@4և���?             ,@2       3       
             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     &@������������������������       �                     @@7       @                    �?�G�z��?             4@8       ?                    �?������?	             .@9       :       
             �?d}h���?             ,@������������������������       �                     "@;       <                    �?���Q��?             @������������������������       �                      @=       >                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @B       �                    �?�`e-��?�            0s@C       \                    �?hy:v�?�            0p@D       K       
             �?���N8�?             E@E       J                 ����?      �?	             0@F       I                    �?���Q��?             @G       H                    b@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     &@L       Y                   �s@�	j*D�?             :@M       V                   �b@z�G�z�?
             4@N       O                    �?      �?             0@������������������������       �                     @P       U                   �`@"pc�
�?             &@Q       R                   @_@����X�?             @������������������������       �                      @S       T                   Pn@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @W       X                    �?      �?             @������������������������       �                      @������������������������       �                      @Z       [                    �F@�q�q�?             @������������������������       �                      @������������������������       �                     @]       �                 `ff@8��?�A�?�             k@^       q                    �?�����H�?�            �i@_       b                    �?d}h���?)             L@`       a                   `U@��
ц��?	             *@������������������������       �                     @������������������������       �                     @c       p                   �e@(L���?             �E@d       m                    `Q@��(\���?             D@e       l       	             �?�}�+r��?             C@f       g                    c@�?�|�?            �B@������������������������       �                     =@h       k                   �U@      �?              @i       j                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?n       o       
             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @r       �                 033@@�+9\J�?a            �b@s       t                    g@�Z]]Y�?V            �`@������������������������       �                    �B@u       �                   �a@,���$�?>            @X@v       }                    �?ܷ��?��?'             M@w       x                   Pc@      �?             0@������������������������       �        	             *@y       z                 ����?�q�q�?             @������������������������       �                     �?{       |                    �I@      �?              @������������������������       �                     �?������������������������       �                     �?~       �                 ��� @���H��?             E@       �                   �i@�ݜ�?            �C@�       �                    Z@      �?             @������������������������       �                      @�       �                 ����?      �?             @�       �                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �       
             �?�FVQ&�?            �@@������������������������       �        	             .@�       �                    @M@�����H�?             2@������������������������       �                     *@�       �                   0r@���Q��?             @�       �                   @`@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �       	             �? ���J��?            �C@������������������������       �                     B@�       �                    �O@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?������?             1@�       �                    �?�q�q�?             (@�       �       
             �?      �?              @������������������������       �                      @������������������������       �                     @�       �                   �_@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     $@�       �                 pff�?r�q��?             H@�       �                    U@      �?             8@������������������������       �                     @�       �                    �?؇���X�?             5@�       �                   �`@�IєX�?
             1@������������������������       �                      @�       �                    �?�����H�?             "@������������������������       �                     @�       �                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                 pff�?      �?             @������������������������       �                      @������������������������       �                      @�       �                   P`@�q�q�?             8@�       �                    �?և���X�?             ,@������������������������       �                     @�       �                 `ff�?�eP*L��?             &@������������������������       �                     @�       �                   �^@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     $@�       �                    �?
�8q���?Z             a@�       �                    �?���N8�?D            @Z@�       �                     R@p�qG�?>             X@�       �                   �b@��s��?=            �W@������������������������       �                    �G@�       �                    �G@�8��8��?             H@������������������������       �                     :@�       �                    �?"pc�
�?             6@������������������������       �                     @�       �                   0c@�}�+r��?             3@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     0@������������������������       �                     �?������������������������       �                     "@�       �                   �^@     ��?             @@������������������������       �                     @�       �                   �n@� �	��?             9@������������������������       �                     "@�       �                   r@     ��?	             0@�       �                    d@8�Z$���?             *@�       �                    �?�8��8��?             (@������������������������       �                     "@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @rM  trN  bh�h"h#K �rO  h%�rP  RrQ  (KK�KK�rR  hZ�B0        s@     �w@      h@     pv@     �`@     �[@     �\@      7@      Z@       @               @      Z@      @     �X@      @     �W@       @      :@             @Q@       @     �J@              0@       @      (@       @      (@                       @      @              @      @      @      @      @                      @      �?              @      �?              �?      @              &@      .@              @      &@      (@               @      &@      @      &@       @      &@      �?      @              @      �?              �?      @                      �?               @      2@      V@      @     �S@      @      @      @               @      @              @       @              �?      S@      �?      F@              ?@      �?      *@      �?       @               @      �?                      &@              @@      &@      "@      &@      @      &@      @      "@               @      @               @       @      �?       @                      �?              �?              @     �M@      o@     �@@     @l@      $@      @@       @      ,@       @      @       @      �?       @                      �?               @              &@       @      2@      @      0@       @      ,@              @       @      "@       @      @               @       @      @       @                      @              @       @       @       @                       @      @       @               @      @              7@     @h@      7@      g@      (@      F@      @      @              @      @              @     �B@      @     �B@       @      B@      �?      B@              =@      �?      @      �?      �?              �?      �?                      @      �?              �?      �?              �?      �?              @              &@     �a@      @     �_@             �B@      @     �V@      @      J@      �?      .@              *@      �?       @              �?      �?      �?              �?      �?              @     �B@      @      A@      @      @       @              �?      @      �?      �?      �?                      �?               @       @      ?@              .@       @      0@              *@       @      @       @      �?              �?       @                       @              @      �?      C@              B@      �?       @      �?                       @      @      *@      @       @       @      @       @                      @       @       @       @                       @              @              $@      :@      6@      2@      @              @      2@      @      0@      �?       @               @      �?      @              �?      �?      �?                      �?       @       @       @                       @       @      0@       @      @      @              @      @              @      @      @              @      @                      $@     �\@      7@      Y@      @     �V@      @     �V@      @     �G@              F@      @      :@              2@      @              @      2@      �?       @      �?              �?       @              0@                      �?      "@              ,@      2@              @      ,@      &@      "@              @      &@       @      &@      �?      &@              "@      �?       @      �?                       @      �?              @        rS  trT  bubhhubh)�rU  }rV  (hhh	h
hNhKhKhG        hh hNhJg}�XhG        hNhG        h@KhAKhBh"h#K �rW  h%�rX  RrY  (KK�rZ  hZ�C              �?r[  tr\  bhNh^hIC       r]  �r^  Rr_  hbKhchdKh"h#K �r`  h%�ra  Rrb  (KK�rc  hI�C       rd  tre  bK�rf  Rrg  }rh  (hKhnK�hoh"h#K �ri  h%�rj  Rrk  (KK�rl  hv�B81         �                    �?z��V���?�           ��@       �                   �b@�y�ʍ+�?b           @�@       l                    �?^����?           �z@                          �_@�j����?�            0v@                        `ff�?P���Q�?=             Y@                        ����?p�C��?7            �V@                          �O@$�q-�?             :@       	                    �?HP�s��?             9@������������������������       �                     4@
                          �X@���Q��?             @������������������������       �                      @                           �L@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �        %            @P@                           �?�q�q�?             "@������������������������       �                      @                           �?և���X�?             @                          @Z@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @       ]                    �?������?�            �o@       T                   pb@|�%�9��?x             i@       -                    �?D�N�dC�?m            �f@       (                    a@��
ц��?             :@                          �`@ҳ�wY;�?             1@������������������������       �                     @       #                   @m@      �?             (@       "       	             �?����X�?             @        !                    �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @$       %                    �?z�G�z�?             @������������������������       �                     @&       '                   `^@      �?              @������������������������       �                     �?������������������������       �                     �?)       ,                   0a@�����H�?             "@*       +       
             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @.       M                   �c@��)�G��?[            �c@/       <                   0j@P���Q�?Q            �a@0       ;                    �?PN��T'�?             ;@1       :                 ����?��s����?             5@2       5                   @_@�q�q�?             (@3       4                   �Z@      �?              @������������������������       �                     �?������������������������       �                     @6       7                   �_@      �?             @������������������������       �                      @8       9                   0g@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@������������������������       �                     @=       H                    �O@ T���v�?=            @\@>       G                   �l@�L��ȕ?4            @W@?       @                    @K@ 7���B�?             ;@������������������������       �                     *@A       B                    �?@4և���?	             ,@������������������������       �                     @C       F                     L@�����H�?             "@D       E                   �k@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �        %            �P@I       J                   (p@ףp=
�?	             4@������������������������       �                     (@K       L                   �p@      �?              @������������������������       �                      @������������������������       �                     @N       O                   �[@      �?
             0@������������������������       �                      @P       S                   Pd@      �?              @Q       R                   �u@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @U       \                   �b@�����?             3@V       [                    �M@�q�q�?             "@W       X                 433�?      �?              @������������������������       �                     @Y       Z                    @      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?������������������������       �                     $@^       _                    �?�E��ӭ�?#             K@������������������������       �                     B@`       g                    �?r�q��?             2@a       f       	             �?؇���X�?	             ,@b       c                   `a@$�q-�?             *@������������������������       �                     $@d       e                   �k@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?h       i                   �p@      �?             @������������������������       �                      @j       k                   `@      �?              @������������������������       �                     �?������������������������       �                     �?m       x                    �?L�qA��?6            �R@n       u                    �?�����?             E@o       r                    �?�L���?            �B@p       q                    �Q@Pa�	�?            �@@������������������������       �                     @@������������������������       �                     �?s       t                    �Q@      �?             @������������������������       �                      @������������������������       �                      @v       w                    ^@z�G�z�?             @������������������������       �                     �?������������������������       �                     @y       �                   �`@���!pc�?            �@@z       �                    �?��
ц��?
             *@{       �                    �?�eP*L��?	             &@|       }                   �Z@�q�q�?             "@������������������������       �                      @~                           �O@؇���X�?             @������������������������       �                     @�       �                 `ff�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                   @]@R���Q�?             4@������������������������       �                     �?�       �                   �m@�KM�]�?             3@������������������������       �        
             (@�       �                   o@����X�?             @������������������������       �                      @������������������������       �                     @�       �                 ���@��6}��?T            �^@�       �                    T@��m��?O            �\@�       �                 ���ܿ����X�?             @������������������������       �                      @������������������������       �                     @�       �                    �?0@�t�?K            �Z@�       �                    �?��]�T��?!            �D@�       �                 @33�?X�<ݚ�?             "@������������������������       �                     @�       �                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                   �g@     ��?             @@������������������������       �                     @�       �       
             �?X�Cc�?             <@�       �                   0j@�q�q�?	             "@������������������������       �                     �?�       �                    �?      �?              @�       �                   `\@؇���X�?             @�       �                   �c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                   l@p�ݯ��?             3@�       �                    @C@      �?              @������������������������       �                     �?�       �                    �?����X�?             @������������������������       �                     �?�       �                    i@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                    �?"pc�
�?	             &@������������������������       �                      @�       �                 ����?�q�q�?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                    �?�U�=���?*            �P@������������������������       �                     �I@�       �                    �?�q�q�?
             .@�       �                    �?      �?             (@�       �       
             �?r�q��?             @������������������������       �                     @�       �                    �F@�q�q�?             @������������������������       �                     �?�       �                   �c@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                     G@�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                   `@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   n@      �?              @������������������������       �                     @������������������������       �                     �?�       �                   `l@0Lj����?V             a@�       �                 ����?���U�?$            �L@�       �                   �P@ �Jj�G�?"            �K@�       �       
             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      J@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?l������?2            �S@�       �                    �?�����H�?'            �O@������������������������       �                     @�       �                    _@����˵�?&            �M@�       �       
             �?      �?             8@������������������������       �                     @�       �                    �?r�q��?             2@������������������������       �                     @�       �                   �^@���!pc�?             &@������������������������       �                      @������������������������       �                     @������������������������       �                    �A@�       �                    �?      �?             0@�       �                   @_@      �?              @������������������������       �                      @������������������������       �                     @������������������������       �                      @rm  trn  bh�h"h#K �ro  h%�rp  Rrq  (KK�KK�rr  hZ�B       pt@     �v@     @j@     `u@      ^@     `s@     @R@     �q@      @     �W@       @     @V@       @      8@       @      7@              4@       @      @               @       @      �?       @                      �?              �?             @P@      @      @               @      @      @      �?      @      �?                      @       @              Q@     `g@      =@     �e@      7@     �c@      (@      ,@      &@      @      @              @      @      @       @      @       @               @      @               @              �?      @              @      �?      �?              �?      �?              �?       @      �?      �?      �?                      �?              @      &@      b@      @     �`@      @      7@      @      1@      @       @      �?      @      �?                      @      @      �?       @              �?      �?      �?                      �?              "@              @      @     �[@      �?      W@      �?      :@              *@      �?      *@              @      �?       @      �?      @              @      �?                      @             �P@       @      2@              (@       @      @       @                      @      @      (@               @      @      @      @      �?      @                      �?              @      @      *@      @      @      @       @      @               @       @               @       @                      �?              $@     �C@      .@      B@              @      .@       @      (@      �?      (@              $@      �?       @      �?                       @      �?              �?      @               @      �?      �?      �?                      �?     �G@      <@      C@      @      A@      @      @@      �?      @@                      �?       @       @               @       @              @      �?              �?      @              "@      8@      @      @      @      @      @      @               @      @      �?      @              �?      �?      �?                      �?               @               @      @      1@      �?               @      1@              (@       @      @       @                      @     �V@      @@     @V@      9@       @      @       @                      @     �U@      4@      :@      .@      @      @              @      @      �?      @                      �?      6@      $@      @              2@      $@      @      @              �?      @       @      @      �?      �?      �?              �?      �?              @                      �?      (@      @      @      @      �?               @      @      �?              �?      @      �?                      @      "@       @       @              �?       @      �?      �?      �?                      �?              �?     �N@      @     �I@              $@      @      "@      @      @      �?      @               @      �?      �?              �?      �?              �?      �?              @       @      @                       @      �?       @      �?                       @      �?      @              @      �?             @]@      3@     �K@       @      K@      �?       @      �?       @                      �?      J@              �?      �?      �?                      �?      O@      1@      L@      @              @      L@      @      5@      @      @              .@      @      @               @      @       @                      @     �A@              @      $@      @       @               @      @                       @rs  trt  bubhhubh)�ru  }rv  (hhh	h
hNhKhKhG        hh hNhJ	�tlhG        hNhG        h@KhAKhBh"h#K �rw  h%�rx  Rry  (KK�rz  hZ�C              �?r{  tr|  bhNh^hIC       r}  �r~  Rr  hbKhchdKh"h#K �r�  h%�r�  Rr�  (KK�r�  hI�C       r�  tr�  bK�r�  Rr�  }r�  (hKhnK�hoh"h#K �r�  h%�r�  Rr�  (KKǅr�  hv�B�+         0                   �d@�#�Ѵ��?�           ��@                           �?��K˱F�?_            �a@                           �?�ګH9�?,            �Q@                           �?`2U0*��?             9@������������������������       �                     8@������������������������       �                     �?                          �c@nM`����?             G@                           `@��V#�?            �E@	                           �I@�㙢�c�?             7@
                           _@���Q��?             $@                          �]@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     *@                          �`@      �?             4@                        033�?r�q��?             @                           P@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                           �?X�Cc�?
             ,@                           I@      �?             $@                        ����?����X�?             @                            B@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @        -                    @�n���?3             R@!       *                   �a@�nkK�?1            @Q@"       #                    �? �.�?Ƞ?,             N@������������������������       �        &             K@$       %                   `]@r�q��?             @������������������������       �                     @&       )                    �?�q�q�?             @'       (                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?+       ,                    �?�<ݚ�?             "@������������������������       �                      @������������������������       �                     @.       /       
             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?1       d                   �`@Lm�&��?T           �@2       ?                    �?��w�r\�?�            `k@3       >       	             �?������?             >@4       9                    `@�	j*D�?             :@5       8                    �?��S�ۿ?             .@6       7                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     (@:       ;                    �?���|���?             &@������������������������       �                     @<       =                   �]@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     @@       O                    �?�YTV��?s            �g@A       B                 ����?j���� �?            �I@������������������������       �                     6@C       H       
             �?�c�Α�?             =@D       G                   �_@؇���X�?             5@E       F       	             �?�z�G��?             $@������������������������       �                     @������������������������       �                     @������������������������       �                     &@I       J                    �?      �?              @������������������������       �                     @K       L                    �M@���Q��?             @������������������������       �                     �?M       N                     R@      �?             @������������������������       �                     @������������������������       �                     �?P       S                    �D@��.N"Ҭ?T            @a@Q       R                   ``@      �?              @������������������������       �                     �?������������������������       �                     �?T       _                 ���@�����?R             a@U       ^                    �?@�n�1�?J            @_@V       W                    �?p� V�?9            �Y@������������������������       �        /            �U@X       Y                   �s@      �?
             0@������������������������       �                     $@Z       [                    �?�q�q�?             @������������������������       �                      @\       ]                   �^@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     6@`       a                    �?�C��2(�?             &@������������������������       �                      @b       c                   p`@�q�q�?             @������������������������       �                     �?������������������������       �                      @e       �                    �?��0�=8�?�            `t@f       �                    �?���H��?�            @j@g       r                   �\@��?}�?w             g@h       q                   @e@@�0�!��?             A@i       n                    �?��+7��?             7@j       k                   �b@�q�q�?             .@������������������������       �                     "@l       m                    �?r�q��?             @������������������������       �                     �?������������������������       �                     @o       p                    @L@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     &@s       t                    �?P-�T6��?c            �b@������������������������       �                    �B@u       v                    d@�}�+r��?L            �\@������������������������       �        )            �M@w       �                    @L@lGts��?#            �K@x                           �?@��8��?             H@y       z                   �^@�g�y��?             ?@������������������������       �        
             .@{       ~                   �j@      �?             0@|       }                   �_@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     (@������������������������       �        
             1@�       �                   0k@����X�?             @�       �                   �i@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �?�q�����?             9@�       �                   �p@
;&����?             7@�       �                 033@�t����?             1@�       �                   @b@؇���X�?	             ,@������������������������       �                     �?�       �                    �I@$�q-�?             *@������������������������       �                     $@�       �                    @K@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                      @�       �                    �?�m�q:@�?C             ]@�       �                    �?�xGZ���?            �A@�       �                    �?8����?             7@�       �                 ����?      �?              @������������������������       �                      @�       �                   @_@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                    �?�r����?
             .@�       �                   �l@8�Z$���?             *@������������������������       �                      @������������������������       �                     &@������������������������       �                      @������������������������       �                     (@�       �                   �f@���R�?/            @T@�       �                   �n@����?-            �S@�       �                    �?8�A�0��?             F@�       �                    �?�'�=z��?            �@@�       �                   �`@      �?
             0@�       �                   �f@      �?              @������������������������       �                     �?�       �                    �?����X�?             @������������������������       �                     �?�       �                   pl@r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                   �j@      �?              @������������������������       �                     @�       �                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    �?�t����?	             1@�       �                   �_@r�q��?             (@�       �                   �^@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                     K@���Q��?             @�       �                   Pj@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                    ^@�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@�       �                   0p@г�wY;�?             A@�       �                   p@ףp=
�?             $@������������������������       �                      @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     8@������������������������       �                     @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KK�KK�r�  hZ�Bp       s@     �w@      7@      ^@      2@     �J@      �?      8@              8@      �?              1@      =@      ,@      =@      @      3@      @      @      �?      @      �?                      @      @                      *@      $@      $@      @      �?      �?      �?              �?      �?              @              @      "@      @      @       @      @       @      �?              �?       @                      @      @                      @      @              @     �P@      @     �P@      �?     �M@              K@      �?      @              @      �?       @      �?      �?      �?                      �?              �?       @      @       @                      @       @      �?       @                      �?     �q@     pp@      L@     `d@      6@       @      2@       @      ,@      �?       @      �?       @                      �?      (@              @      @      @              �?      @              @      �?              @              A@     `c@      >@      5@      6@               @      5@      @      2@      @      @              @      @                      &@      @      @      @               @      @      �?              �?      @              @      �?              @     �`@      �?      �?              �?      �?              @     �`@       @     �^@       @     @Y@             �U@       @      ,@              $@       @      @               @       @       @       @                       @              6@      �?      $@               @      �?       @      �?                       @     @l@      Y@      g@      9@     �e@      (@      <@      @      1@      @      $@      @      "@              �?      @      �?                      @      @      �?      @                      �?      &@              b@      @     �B@              [@      @     �M@             �H@      @     �G@      �?      >@      �?      .@              .@      �?      @      �?              �?      @              (@              1@               @      @       @      �?              �?       @                      @      (@      *@      (@      &@      (@      @      (@       @              �?      (@      �?      $@               @      �?              �?       @                      @              @               @     �D@     �R@      3@      0@      @      0@      @      @               @      @      �?              �?      @               @      *@       @      &@       @                      &@               @      (@              6@     �M@      3@     �M@      2@      :@      1@      0@      (@      @      @      @              �?      @       @              �?      @      �?      @                      �?      @      �?      @              @      �?      @                      �?      @      (@       @      $@       @      @              @       @                      @      @       @      �?       @               @      �?               @              �?      $@      �?                      $@      �?     �@@      �?      "@               @      �?      �?      �?                      �?              8@      @        r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ�ޡhG        hNhG        h@KhAKhBh"h#K �r�  h%�r�  Rr�  (KK�r�  hZ�C              �?r�  tr�  bhNh^hIC       r�  �r�  Rr�  hbKhchdKh"h#K �r�  h%�r�  Rr�  (KK�r�  hI�C       r�  tr�  bK�r�  Rr�  }r�  (hKhnMhoh"h#K �r�  h%�r�  Rr�  (KM�r�  hv�B�:         �                    �?�H��3��?�           ��@       o                    �?0}&Ν>�?           �x@       `                    �?�L"��?�            t@       G                    �L@�X�3�m�?�            pr@                           �?�W��}�?c            �c@                           �?П[;U��?             =@������������������������       �                     �?                          w@���>4��?             <@	              	             �?8�A�0��?             6@
                          Pb@�G�z��?             4@                           b@ҳ�wY;�?	             1@                        ����?      �?              @������������������������       �                     @������������������������       �                     @              
             �?�<ݚ�?             "@                        ��� @z�G�z�?             @������������������������       �                     @������������������������       �                     �?                          `\@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                     @                          �U@�?�<��?T            @`@������������������������       �                      @       B                    �?     ��?S             `@       =       	             �?(L���?:            �U@                           �?      �?4             T@������������������������       �                      @                           �Z@4?,R��?/             R@������������������������       �                     �?!       *                    �?��UV�?.            �Q@"       #                 ����?������?             1@������������������������       �                     $@$       %       
             �?և���X�?             @������������������������       �                     �?&       '                   �^@�q�q�?             @������������������������       �                     �?(       )                 ����?z�G�z�?             @������������������������       �                     @������������������������       �                     �?+       0                   �f@h�WH��?#             K@,       -                   @_@      �?             (@������������������������       �                     @.       /                    �?      �?             @������������������������       �                     @������������������������       �                     @1       2                    @J@���N8�?             E@������������������������       �                     >@3       :                    @r�q��?	             (@4       9                    �?ףp=
�?             $@5       6                   @[@z�G�z�?             @������������������������       �                     @7       8                     K@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @;       <                   p@      �?              @������������������������       �                     �?������������������������       �                     �?>       A       
             �?�q�q�?             @?       @                    @I@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @C       D                    r@���N8�?             E@������������������������       �                     >@E       F                    �?r�q��?             (@������������������������       �                      @������������������������       �                     $@H       U                   �b@�wY;��?Z             a@I       J                 033�?�]0��<�?P            �^@������������������������       �        2            �Q@K       P                    �?�:�]��?            �I@L       M                   �b@؇���X�?
             ,@������������������������       �                     "@N       O                     P@���Q��?             @������������������������       �                     @������������������������       �                      @Q       R                   Hr@@-�_ .�?            �B@������������������������       �                    �@@S       T       
             �?      �?             @������������������������       �                      @������������������������       �                      @V       _                    �?d}h���?
             ,@W       X                    ]@      �?             @������������������������       �                      @Y       ^       
             �?      �?             @Z       [                   pp@�q�q�?             @������������������������       �                     �?\       ]                   d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @a       h                    n@
j*D>�?             :@b       e                    �?d}h���?
             ,@c       d                   �[@�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@f       g                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @i       n                 ����?�q�q�?             (@j       m                    �?X�<ݚ�?             "@k       l                    �?      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     @p       s                    @G@��J�fj�?2            �R@q       r                   @b@�C��2(�?	             &@������������������������       �                     $@������������������������       �                     �?t       {                    �?b����?)            �O@u       z                   @b@�<ݚ�?             "@v       y                    �?�q�q�?             @w       x                 ����?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @|       �                   �d@�E��ӭ�?"             K@}       �                    �?      �?!             J@~                           �J@x�����?            �C@������������������������       �                     &@�       �                    �?����X�?             <@�       �                 `ff�?�LQ�1	�?             7@�       �                    �?���|���?             &@�       �                    @L@r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                     N@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                    �N@�8��8��?             (@������������������������       �                     @�       �                    �?z�G�z�?             @������������������������       �                      @�       �                   Pa@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   Pj@�n_Y�K�?	             *@�       �                    �M@r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                   �^@և���X�?             @������������������������       �                     @�       �                    �P@      �?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                    �K@Z��G{R�?�            Pr@�       �                    �?|�5�L�?�            �k@�       �                 033�? �M*k�?�            �h@�       �                 833�?�+?�?�            �g@�       �                    P@�&=�w��?n            �c@�       �       
             �?      �?             @�       �                    @D@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                    @F@ ���l��?k            `c@�       �                    �E@��`qM|�?;            �T@�       �                    �C@������?3             R@������������������������       �                    �D@�       �       
             �?`Jj��?             ?@�       �                    \@z�G�z�?             @�       �                   �b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    @D@ ��WV�?             :@�       �                   f@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     7@�       �                   �i@"pc�
�?             &@������������������������       �                     �?�       �                    �?ףp=
�?             $@�       �                    �?      �?              @�       �                   Hq@؇���X�?             @������������������������       �                     @�       �       
             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �        0             R@�       �                    �?�חF�P�?             ?@������������������������       �                      @�       �                    �?��<b���?             7@�       �                    �?�t����?
             1@�       �                 hff�?      �?             $@������������������������       �                      @�       �                     I@      �?              @������������������������       �                      @�       �                   �`@r�q��?             @�       �                   `]@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �       	             �?����X�?             @�       �                    ^@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�       �                    I@\X��t�?             7@������������������������       �                     $@�       �                   �s@�θ�?             *@�       �       
             �?r�q��?
             (@������������������������       �                     @�       �                    �?�<ݚ�?             "@�       �                 033�?����X�?             @�       �                 `ff�?z�G�z�?             @�       �                   @]@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�                          �?P�t��?0            @R@�                          `R@�c�����?"            �J@�       �                    g@��[�8��?!            �I@�       �       
             �?X�<ݚ�?             "@������������������������       �                     @�       �                     P@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    �?r�q��?             E@�       �                   0d@�C��2(�?            �@@�       �                    �? 7���B�?             ;@������������������������       �                     7@�       �                    q@      �?             @�       �                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    �?�q�q�?             @�       �                   @e@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �                   �_@X�<ݚ�?             "@������������������������       �                     @�                          �`@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @                        �V@z�G�z�?             4@������������������������       �                     (@                         �L@      �?              @������������������������       �                      @                         `P@�q�q�?             @      	                  �`@z�G�z�?             @������������������������       �                      @
                         �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KMKK�r�  hZ�B�       �s@      w@     �T@     �s@     �I@     �p@      B@     0p@      =@     @`@      *@      0@              �?      *@      .@      *@      "@      &@      "@      &@      @      @      @      @                      @      @       @      @      �?      @                      �?      @      �?              �?      @                      @       @                      @      0@     �\@       @              ,@     �\@      (@     �R@      $@     �Q@               @      $@      O@      �?              "@      O@      @      *@              $@      @      @              �?      @       @              �?      @      �?      @                      �?      @     �H@      @      "@              @      @      @              @      @               @      D@              >@       @      $@      �?      "@      �?      @              @      �?      �?              �?      �?                      @      �?      �?              �?      �?               @      @       @       @               @       @                       @       @      D@              >@       @      $@       @                      $@      @      `@      @     �]@             �Q@      @     �G@       @      (@              "@       @      @              @       @               @     �A@             �@@       @       @               @       @              @      &@      @      @               @      @      �?       @      �?      �?              �?      �?      �?                      �?      �?                       @      .@      &@      &@      @      $@      �?              �?      $@              �?       @      �?                       @      @       @      @      @      @      @      @                      @              �?              @      @@      E@      $@      �?      $@                      �?      6@     �D@      @       @      �?       @      �?      �?              �?      �?                      �?      @              .@     �C@      *@     �C@       @      ?@              &@       @      4@       @      .@      @      @      @      �?      @                      �?       @      @       @                      @      �?      &@              @      �?      @               @      �?       @               @      �?                      @      @       @      �?      @              @      �?              @      @      @              �?      @      �?      �?      �?                      �?               @       @             `m@      M@     �g@      =@     �f@      0@     `f@      &@      c@      @       @       @      �?       @               @      �?              �?             �b@      @     �S@      @     �Q@       @     �D@              =@       @      @      �?      �?      �?      �?                      �?      @              9@      �?       @      �?       @                      �?      7@              "@       @              �?      "@      �?      @      �?      @      �?      @              �?      �?              �?      �?              �?               @              R@              :@      @       @              2@      @      (@      @      @      @               @      @      @               @      @      �?      �?      �?      �?                      �?      @              @              @               @      @      �?      @              @      �?              �?              $@      *@              $@      $@      @      $@       @      @              @       @      @       @      @      �?      @      �?      @                      �?      �?              �?      �?      �?                      �?       @                      �?      F@      =@      D@      *@      D@      &@      @      @      @              �?      @              @      �?             �A@      @      >@      @      :@      �?      7@              @      �?      �?      �?              �?      �?               @              @       @      @       @               @      @              �?              @      @      @               @      @              @       @                       @      @      0@              (@      @      @       @               @      @      �?      @               @      �?       @               @      �?              �?        r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJQY%hG        hNhG        h@KhAKhBh"h#K �r�  h%�r�  Rr�  (KK�r�  hZ�C              �?r�  tr�  bhNh^hIC       r�  �r�  Rr�  hbKhchdKh"h#K �r�  h%�r�  Rr�  (KK�r�  hI�C       r�  tr�  bK�r�  Rr�  }r�  (hKhnK�hoh"h#K �r�  h%�r�  Rr�  (KKхr�  hv�B�-         �                   �a@L��&�?�           ��@       K                    �?d�����?D           �@                           �?l��q �?�            Pp@                          �m@�<ݚ�?             B@                           �?�>����?             ;@                           U@      �?             0@                          @\@����X�?             @������������������������       �                      @	       
                   �V@���Q��?             @������������������������       �                     �?                           �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     "@������������������������       �                     &@                          �^@�q�q�?             "@������������������������       �                      @                          �`@؇���X�?             @������������������������       �                     @������������������������       �                     �?       <                    �?
�O3���?�             l@       ;                    �R@T�\�9�?y             g@                           I@x93c�?x            �f@                           �?�q�q�?	             (@                          �d@      �?              @������������������������       �                     @������������������������       �                      @                           �?      �?             @������������������������       �                      @������������������������       �                      @       *                    �I@���U�?o            `e@        )                   �[@@�n���?A            �Y@!       "                    �? ��WV�?             :@������������������������       �        	             0@#       (                    �?ףp=
�?             $@$       %                   �c@�����H�?             "@������������������������       �                     @&       '                   �j@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �        1            @S@+       0                    @J@����p�?.             Q@,       /                   �d@d}h���?             ,@-       .                   Pc@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     @1       6                   �? 7���B�?'             K@2       3                   xs@����?�?!            �F@������������������������       �                     D@4       5                    `@z�G�z�?             @������������������������       �                     @������������������������       �                     �?7       8                    �?�����H�?             "@������������������������       �                     @9       :                   d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @=       >                   �_@      �?             D@������������������������       �                     1@?       @                    �?\X��t�?             7@������������������������       �                     @A       J                    �?�����?             3@B       E                   �`@     ��?             0@C       D                   �r@�q�q�?             @������������������������       �                      @������������������������       �                     �?F       G                    �?$�q-�?	             *@������������������������       �                     $@H       I                    �G@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @L       q       
             �?w�=B�?�            �o@M       T                    �?\��<�|�?=            �W@N       S                    �?�q�q�?	             (@O       R                   �b@z�G�z�?             $@P       Q                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                      @U       \                   �?b:�&���?4            �T@V       [                   �?և���X�?             ,@W       Z                    �?z�G�z�?             $@X       Y                    ^@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     @]       l                   �c@�LQ�1	�?,            @Q@^       _                   �i@ ,��-�?$            �M@������������������������       �                     ;@`       a                    �?      �?             @@������������������������       �        
             1@b       k                    @������?             .@c       d                    �H@d}h���?
             ,@������������������������       �                      @e       j                    �?�8��8��?	             (@f       i                   �`@ףp=
�?             $@g       h                   �l@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                     �?m       n                    �L@      �?             $@������������������������       �                     @o       p                   �\@r�q��?             @������������������������       �                     �?������������������������       �                     @r       s                   �c@Ld����?^            �c@������������������������       �                    �I@t       �                    �?�#ʆA��??            �Z@u       v                   pl@��.k���?             1@������������������������       �                     @w       |                    �H@�q�q�?             (@x       {                    �?���Q��?             @y       z                   �n@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?}       ~                 433�?؇���X�?             @������������������������       �                     @       �                 ����?      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �?��~l�?3            @V@�       �                 ����?|��"J�?.            @T@�       �                 ����?J�8���?             =@������������������������       �        
             3@������������������������       �                     $@�       �                   ``@ȵHPS!�?!             J@�       �                    �?�MI8d�?            �B@�       �                   Xr@      �?             @@������������������������       �                     :@�       �                    @I@�q�q�?             @�       �                   @_@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �O@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     .@�       �                     @      �?              @�       �                 ����?r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                    �?���<��?r            �e@�       �                    �?`�Q��?R            @_@�       �                    �?���W���?5            �U@�       �       	             �?�+$�jP�?             ;@�       �       
             �?�LQ�1	�?             7@�       �                 ����?�θ�?             *@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     "@������������������������       �                     $@�       �                    �P@      �?             @������������������������       �                      @������������������������       �                      @�       �                    �? ,��-�?(            �M@�       �                    �H@��<b�ƥ?!             G@�       �                   Pl@؇���X�?             @������������������������       �                     @�       �                   �p@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                    �C@�       �                 ����?�θ�?             *@�       �                    �M@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @�       �                 ����?x�����?            �C@�       �       	             �?r�q��?             B@�       �                   Pc@�n`���?             ?@�       �                    �?X�Cc�?
             ,@�       �                   �m@X�<ݚ�?             "@������������������������       �                     @�       �                   �p@z�G�z�?             @������������������������       �                      @�       �                 ����?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �O@�IєX�?             1@�       �                   `X@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     $@������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?H%u��?              I@�       �                    �?����?�?            �F@�       �       	             �?�nkK�?             7@������������������������       �                     5@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     6@������������������������       �                     @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KK�KK�r�  hZ�B       �q@      y@      n@     q@     `g@     �R@       @      <@       @      9@       @      ,@       @      @               @       @      @      �?              �?      @              @      �?                      "@              &@      @      @               @      @      �?      @                      �?     `f@      G@      e@      0@      e@      ,@      @       @       @      @              @       @               @       @       @                       @     �d@      @     �Y@      �?      9@      �?      0@              "@      �?       @      �?      @              �?      �?              �?      �?              �?             @S@             �O@      @      &@      @      @      @      @                      @      @              J@       @      F@      �?      D@              @      �?      @                      �?       @      �?      @              �?      �?              �?      �?                       @      $@      >@              1@      $@      *@      @              @      *@      @      *@       @      �?       @                      �?      �?      (@              $@      �?       @      �?                       @      @             �J@     �h@      7@      R@       @      @       @       @       @       @       @                       @      @                       @      .@      Q@      @       @       @       @       @       @       @                       @              @      @              "@      N@      @     �K@              ;@      @      <@              1@      @      &@      @      &@       @              �?      &@      �?      "@      �?      @      �?                      @              @               @      �?              @      @      @              �?      @      �?                      @      >@     �_@             �I@      >@      S@      "@       @      @              @       @      @       @       @       @       @                       @      �?              �?      @              @      �?      @      �?                      @      5@      Q@      0@     @P@      $@      3@              3@      $@              @      G@      @      ?@       @      >@              :@       @      @       @      �?              �?       @                      @      @      �?      @                      �?              .@      @      @      @      �?              �?      @                       @      G@      `@      D@     @U@      "@     @S@      @      6@      @      4@      @      $@      @      �?      @                      �?              "@              $@       @       @       @                       @      @     �K@      �?     �F@      �?      @              @      �?      @      �?                      @             �C@      @      $@      @       @      @                       @               @      ?@       @      >@      @      9@      @      "@      @      @      @              @      @      �?       @               @      �?              �?       @              @              0@      �?      @      �?              �?      @              $@              @              �?       @      �?                       @      @      F@      �?      F@      �?      6@              5@      �?      �?      �?                      �?              6@      @        r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ��fbhG        hNhG        h@KhAKhBh"h#K �r�  h%�r�  Rr�  (KK�r�  hZ�C              �?r�  tr�  bhNh^hIC       r�  �r�  Rr�  hbKhchdKh"h#K �r�  h%�r�  Rr�  (KK�r�  hI�C       r�  tr�  bK�r�  Rr�  }r�  (hKhnK�hoh"h#K �r�  h%�r�  Rr�  (KK݅r�  hv�BX0                             _@�կZ���?�           ��@                          P`@�U�=���?R            �`@                           �?@��,B�?9            �V@                          `X@ ���J��?            �C@                           �?؇���X�?             @������������������������       �                      @       
                    �?z�G�z�?             @       	                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @@������������������������       �        "             J@                           �?��P���?            �D@                           c@�q�q�?             2@                           �?؇���X�?
             ,@              
             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     &@������������������������       �                     @                          �c@�LQ�1	�?             7@������������������������       �        
             1@              
             �?      �?             @                          0d@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?       >                    �?�W���?b           `�@       )                    �?b���f�?W             a@       "                   Pe@�d���?7            �U@        !       
             �?      �?              @������������������������       �                     �?������������������������       �                     �?#       $                   �`@`��>�ϗ?5            @U@������������������������       �                     H@%       &                   �s@�?�|�?            �B@������������������������       �                     @@'       (                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?*       =                    �?z�):���?              I@+       <                    `P@X�Cc�?             E@,       1                    �?և���X�?            �A@-       0                    �?z�G�z�?             4@.       /                   �a@������?             1@������������������������       �                     *@������������������������       �                     @������������������������       �                     @2       3       
             �?������?	             .@������������������������       �                     @4       7                   �`@�q�q�?             (@5       6                    @E@      �?             @������������������������       �                     �?������������������������       �                     @8       9                 433�?      �?              @������������������������       �                     @:       ;                   �k@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @?       �                    �K@��f帩�?           0z@@       {                    �?�>4ևF�?�             l@A       r                    �?$���'w�?c            �a@B       q                    @J@�՘���?C            �W@C       p                   h}@0,Tg��?;             U@D       E                     C@R���Q�?:             T@������������������������       �                     $@F       O                    @D@��R[s�?4            �Q@G       J                    m@�eP*L��?             &@H       I                   @`@z�G�z�?             @������������������������       �                     �?������������������������       �                     @K       L                   �b@r�q��?             @������������������������       �                     @M       N                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?P       U                   @`@��$�4��?,            �M@Q       T                   �d@�q�q�?             @R       S                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?V       e                    �?�iʫ{�?'            �J@W       `       
             �?�q��/��?              G@X       _                    �?�q�q�?             (@Y       Z                   0j@և���X�?             @������������������������       �                     @[       ^                 ����?      �?             @\       ]                     G@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @a       b                   �d@г�wY;�?             A@������������������������       �                     7@c       d                    e@�C��2(�?	             &@������������������������       �                     �?������������������������       �                     $@f       g                   �\@և���X�?             @������������������������       �                     �?h       o                   �i@      �?             @i       n                    �?      �?             @j       k                   �a@�q�q�?             @������������������������       �                     �?l       m                   �]@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     &@s       z                    �?      �?              H@t       u                   Pa@�θ�?	             *@������������������������       �                     �?v       y                   �m@r�q��?             (@w       x                   �d@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     "@������������������������       �                    �A@|       �                    �?ڤ���?3            @T@}       ~                    �?���Q��?             4@������������������������       �                     �?       �                   `d@p�ݯ��?
             3@�       �                    �?��
ц��?             *@�       �                   �`@�q�q�?             "@�       �       
             �?      �?             @������������������������       �                     �?�       �                    n@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                 ����?(��+�?(            �N@�       �                   �[@tk~X��?             B@�       �                    b@և���X�?             @������������������������       �                     @������������������������       �                     @�       �                    _@ܷ��?��?             =@�       �                    �?      �?              @�       �                   Pa@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�       �                   �_@���N8�?             5@������������������������       �                     (@�       �                    �E@�����H�?             "@������������������������       �                     �?������������������������       �                      @�       �       
             �?`2U0*��?             9@�       �                    b@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     2@�       �                    �M@��Sݭg�?u            `h@�       �                    �?^�JB=�?0            @T@�       �                    �?     ��?$             P@�       �                    @M@�LQ�1	�?             G@�       �                   �h@��?^�k�?            �A@������������������������       �                     �?������������������������       �                     A@�       �       
             �?�eP*L��?             &@������������������������       �                     �?�       �                   �]@      �?             $@������������������������       �                      @�       �                   �^@      �?              @������������������������       �                     @�       �                   �`@���Q��?             @������������������������       �                     @������������������������       �                      @�       �                   Pk@�<ݚ�?             2@�       �       	             �?$�q-�?             *@������������������������       �                     (@������������������������       �                     �?�       �                    b@���Q��?             @�       �                    �?�q�q�?             @�       �                   ``@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                   Hp@ҳ�wY;�?             1@�       �                   `b@8�Z$���?	             *@�       �                 hff�?�8��8��?             (@������������������������       �                     $@�       �                   @`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �`@r�q��?E            �\@�       �                 ����?�5��
J�?             G@�       �                   �s@���!pc�?             &@�       �                    �?�����H�?             "@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                   �_@�#-���?            �A@������������������������       �                     7@�       �                   @n@      �?	             (@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    �?�t����?*             Q@�       �                    �?���Q��?             4@�       �                    �?      �?              @�       �       	             �?����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �                    �R@r�q��?             (@������������������������       �                     $@������������������������       �                      @������������������������       �                     H@r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KK�KK�r�  hZ�B�       `s@     �w@      $@     �^@      �?     �V@      �?      C@      �?      @               @      �?      @      �?       @               @      �?                       @              @@              J@      "@      @@      @      (@       @      (@       @      �?              �?       @                      &@      @              @      4@              1@      @      @      @       @      @                       @              �?     �r@      p@      \@      9@     @U@       @      �?      �?              �?      �?              U@      �?      H@              B@      �?      @@              @      �?      @                      �?      ;@      7@      ;@      .@      4@      .@      0@      @      *@      @      *@                      @      @              @      &@              @      @       @      @      �?              �?      @              �?      @              @      �?      �?              �?      �?              @                       @     �g@     �l@     @a@     �U@     �]@      9@     @R@      6@      O@      6@      O@      2@      $@              J@      2@      @      @      �?      @      �?                      @      @      �?      @               @      �?       @                      �?      G@      *@       @      @      �?      @              @      �?              �?              F@      "@     �D@      @       @      @      @      @              @      @      �?      �?      �?              �?      �?               @              @             �@@      �?      7@              $@      �?              �?      $@              @      @              �?      @      @      @      �?       @      �?      �?              �?      �?      �?                      �?      �?                       @              @      &@             �F@      @      $@      @              �?      $@       @      �?       @               @      �?              "@             �A@              4@     �N@      (@       @              �?      (@      @      @      @      @      @      �?      @              �?      �?       @      �?                       @      @                      @      @               @     �J@      @      =@      @      @      @                      @      @      :@       @      @      �?      @              @      �?              �?              �?      4@              (@      �?       @      �?                       @      �?      8@      �?      @              @      �?                      2@      I@      b@      ?@      I@      4@      F@      @      D@      �?      A@      �?                      A@      @      @              �?      @      @               @      @      @      @               @      @              @       @              ,@      @      (@      �?      (@                      �?       @      @       @      �?      �?      �?      �?                      �?      �?                       @      &@      @      &@       @      &@      �?      $@              �?      �?      �?                      �?              �?              @      3@     �W@      &@     �A@       @      @       @      �?      @      �?      @                      �?      @                       @      @      @@              7@      @      "@      @      @      @                      @              @       @      N@       @      (@      @       @      @       @               @      @              �?               @      $@              $@       @                      H@r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ$�phG        hNhG        h@KhAKhBh"h#K �r�  h%�r�  Rr�  (KK�r�  hZ�C              �?r�  tr�  bhNh^hIC       r�  �r�  Rr�  hbKhchdKh"h#K �r   h%�r  Rr  (KK�r  hI�C       r  tr  bK�r  Rr  }r  (hKhnK�hoh"h#K �r	  h%�r
  Rr  (KK�r  hv�B�1         R                 ����?v ��?�           ��@       3                    �?�R�[��?�            �t@                            @L@=�J�C�?�            �m@                          �f@�+?�?m            �g@       
                    I@`2U0*��?e            �e@       	                    _@      �?              @                          �d@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @                          �b@ d��?`            �d@������������������������       �        .             T@                           �?`��F:u�?2            �U@                          �\@(�5�f��?-            �S@                          �Z@���!pc�?	             &@������������������������       �                     @                           �G@և���X�?             @                           @E@���Q��?             @              
             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �        $             Q@                           �?      �?              @              
             �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @                          �a@������?             .@������������������������       �                     &@������������������������       �                     @!       2                    �? \� ���?            �H@"       #                   `Q@�����?             C@������������������������       �                     @$       1                    �?������?             A@%       ,                   �b@�LQ�1	�?             7@&       '                   @a@$�q-�?
             *@������������������������       �                     @(       )                   �o@r�q��?             @������������������������       �                     @*       +                    q@�q�q�?             @������������������������       �                     �?������������������������       �                      @-       .                    c@�z�G��?             $@������������������������       �                     @/       0                    �?և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     &@������������������������       �                     &@4       =                    �?�<ݚ�?8            �V@5       6                    �?j���� �?             1@������������������������       �                     @7       8                   b@�θ�?             *@������������������������       �                      @9       :                   �n@�C��2(�?             &@������������������������       �                     @;       <                   pp@      �?             @������������������������       �                     �?������������������������       �                     @>       O                    �?d1<+�C�?-            @R@?       N                   �f@ДX��?*             Q@@       A                    �J@�U�=���?)            �P@������������������������       �                     9@B       E                    �K@,���i�?            �D@C       D                    �?      �?             @������������������������       �                      @������������������������       �                      @F       G                   �f@�L���?            �B@������������������������       �                     9@H       M                    b@      �?	             (@I       L                    @O@և���X�?             @J       K                   Pj@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                      @P       Q                   `\@���Q��?             @������������������������       �                      @������������������������       �                     @S       �                    �?$nW-��?�            pv@T       �                    �?�S����?�            �q@U       �                   �a@����[��?8            �S@V       u                   �b@���Q��?,             N@W       Z                    �?�^�����?            �E@X       Y                   @_@�q�q�?             @������������������������       �                     @������������������������       �                      @[       r                   �`@V������?            �B@\       g                   �p@X�Cc�?             <@]       `                    �?������?             1@^       _                   �o@���Q��?             @������������������������       �                     @������������������������       �                      @a       b       
             �?�8��8��?             (@������������������������       �                     @c       d                   @_@�����H�?             "@������������������������       �                     @e       f                 033@      �?              @������������������������       �                     �?������������������������       �                     �?h       m                   �\@�eP*L��?             &@i       l                   �s@      �?             @j       k                   @_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @n       o                    �?����X�?             @������������������������       �                     @p       q                    �K@      �?             @������������������������       �                      @������������������������       �                      @s       t                   `^@�����H�?             "@������������������������       �                     �?������������������������       �                      @v       w                    @C@ҳ�wY;�?             1@������������������������       �                     �?x       y                    ]@     ��?             0@������������������������       �                     @z       {                   �?8�Z$���?
             *@������������������������       �                     @|                        `ff�?����X�?             @}       ~                   �c@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                 `ff@�X�<ݺ?             2@������������������������       �                     1@������������������������       �                     �?�       �                    �?�Q�1X�?y            �i@�       �                    �?0�,��?j            �f@�       �                    �?�<ݚ�?
             2@�       �                   �`@���|���?             &@�       �                    �I@z�G�z�?             @�       �                   �_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                   �U@�ۊ�̴?`            �d@������������������������       �                     �?�       �                   @i@Ћ����?_            �d@�       �                   `c@     p�?$             P@�       �                    �?Hn�.P��?#             O@�       �                    �?����˵�?"            �M@�       �       
             �?=QcG��?            �G@������������������������       �                     &@�       �                   �h@�8��8��?             B@�       �                   @e@Pa�	�?            �@@������������������������       �                     9@�       �                 `ff @      �?              @�       �                   @`@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     (@������������������������       �                     @������������������������       �                      @�       �                   pa@ �ׁsF�?;             Y@������������������������       �        $             O@�       �                    �?P�Lt�<�?             C@�       �       
             �?���7�?             6@������������������������       �                     @�       �                   �a@�X�<ݺ?             2@�       �                     J@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     &@������������������������       �        	             0@�       �                    �?      �?             8@�       �                   P`@�q�q�?	             (@�       �                    �N@�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                   �a@r�q��?             @������������������������       �                     @�       �                    @G@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    @M@�q�q�?             (@������������������������       �                     @�       �                    �P@�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                    �?(ǯt��?/            �R@�       �       	             �?�2�o�U�?#            �K@�       �                    �?���Q �?             �H@�       �                    �?�s��:��?             C@������������������������       �                     $@�       �                   `b@��>4և�?             <@�       �                    �?8����?             7@�       �                   �n@@�0�!��?             1@�       �                    �?      �?              @�       �                    �?      �?             @�       �                   �`@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     "@�       �                   �d@�q�q�?             @�       �                    _@z�G�z�?             @�       �                   �\@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �       
             �?z�G�z�?             @�       �                   `c@      �?             @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@������������������������       �                     @�       �                    �?�}�+r��?             3@������������������������       �                     �?������������������������       �                     2@r  tr  bh�h"h#K �r  h%�r  Rr  (KK�KK�r  hZ�B0        t@      w@     �m@     @W@      k@      7@     `f@      &@      e@      @      @      @       @      @              @       @              @             `d@      @      T@             �T@      @      S@      @       @      @      @              @      @       @      @       @      �?              �?       @                       @       @              Q@              @      �?      @      �?              �?      @              @              &@      @      &@                      @     �B@      (@      :@      (@              @      :@       @      .@       @      (@      �?      @              @      �?      @               @      �?              �?       @              @      @              @      @      @      @                      @      &@              &@              4@     �Q@      $@      @              @      $@      @               @      $@      �?      @              @      �?              �?      @              $@     �O@      @     �N@      @     �N@              9@      @      B@       @       @               @       @              @      A@              9@      @      "@      @      @      �?      @      �?                      @       @                      @       @              @       @               @      @              U@     0q@     �F@      n@      9@     �J@      8@      B@      *@      >@       @      @              @       @              &@      :@      $@      2@      @      *@      @       @      @                       @      �?      &@              @      �?       @              @      �?      �?      �?                      �?      @      @      �?      @      �?      �?              �?      �?                       @      @       @      @               @       @       @                       @      �?       @      �?                       @      &@      @              �?      &@      @              @      &@       @      @              @       @      �?       @      �?                       @      @              �?      1@              1@      �?              4@     `g@      &@     �e@      @      ,@      @      @      @      �?      �?      �?      �?                      �?      @                      @              @      @     �c@      �?              @     �c@      @     �M@      @     �M@      @      L@      @      F@              &@      @     �@@      �?      @@              9@      �?      @      �?      @              @      �?                      @       @      �?       @                      �?              (@              @       @              �?     �X@              O@      �?     �B@      �?      5@              @      �?      1@      �?      @              @      �?                      &@              0@      "@      .@      @      @      @       @      @                       @      �?      @              @      �?       @      �?                       @      @       @              @      @       @      @                       @     �C@     �A@      C@      1@      @@      1@      5@      1@      $@              &@      1@      @      0@      @      ,@      @      @      @      @      �?       @               @      �?               @      �?              �?       @                       @              "@      @       @      @      �?      �?      �?      �?                      �?      @                      �?      @      �?      @      �?       @      �?       @                      �?      �?              �?              &@              @              �?      2@      �?                      2@r  tr  bubhhubh)�r  }r  (hhh	h
hNhKhKhG        hh hNhJW:+LhG        hNhG        h@KhAKhBh"h#K �r  h%�r  Rr  (KK�r  hZ�C              �?r  tr  bhNh^hIC       r  �r  Rr  hbKhchdKh"h#K �r   h%�r!  Rr"  (KK�r#  hI�C       r$  tr%  bK�r&  Rr'  }r(  (hKhnK�hoh"h#K �r)  h%�r*  Rr+  (KKǅr,  hv�B�+         h                 033�?xa@����?�           ��@       O                    �?�u�ea��?�            �w@                          �\@>��C��?�            �r@                           �?և���X�?             <@������������������������       �        	             (@������������������������       �                     0@                           �?��܂O�?�            q@                          �c@Dc}h��?#             L@	              
             �?���7�?             6@
                        `ff�?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �        
             1@                          �d@��.k���?             A@                          �b@�q�q�?             8@                           �?r�q��?             @������������������������       �                     @                           a@      �?              @������������������������       �                     �?������������������������       �                     �?                           �?r�q��?	             2@                          �c@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     *@                           �D@z�G�z�?             $@������������������������       �                     �?                          �n@�����H�?             "@������������������������       �                      @������������������������       �                     �?       (                    @A@�
���x�?�             k@        %       	             �?�θ�?	             *@!       $                   �c@ףp=
�?             $@"       #       
             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @&       '                 `ff�?�q�q�?             @������������������������       �                     �?������������������������       �                      @)       0                    �?�IєX�?�            �i@*       +                    �L@�J�T�?,            �Q@������������������������       �        "             M@,       /                    �N@8�Z$���?
             *@-       .                   Pe@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     $@1       H                    �?`�bV��?T            �`@2       3                   �h@ą%�E�?7            @V@������������������������       �                     8@4       5                   �h@��ɉ�?*            @P@������������������������       �                     @6       G                    �?��a�n`�?)             O@7       D                    @L@���C��?"            �J@8       C                    �?���.�6�?             G@9       B                   �b@��2(&�?             6@:       A       
             �?�����?             5@;       @       	             �?r�q��?             (@<       =                   Pb@�<ݚ�?             "@������������������������       �                     @>       ?                    e@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     "@������������������������       �                     �?������������������������       �                     8@E       F                    �L@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     "@I       N                   �]@`���i��?             F@J       K                   �R@�����H�?             "@������������������������       �                     @L       M                 pff�?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                    �A@P       U                    �?&:~�Q�?.             S@Q       R                    l@P���Q�?             D@������������������������       �                     8@S       T                 833�?      �?
             0@������������������������       �                     ,@������������������������       �                      @V       Y                   �Z@<ݚ)�?             B@W       X                    ^@      �?             @������������������������       �                     �?������������������������       �                     @Z       _                   `c@      �?             @@[       \                 ����?�IєX�?             1@������������������������       �                     &@]       ^                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?`       a                    �?��S���?	             .@������������������������       �                     @b       g                    �?�q�q�?             (@c       d                   @`@�eP*L��?             &@������������������������       �                     @e       f                   pd@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?i       �                    �?Σq���?�            ps@j       �                   �b@T��o��?�            Pp@k       l                   Pe@ �Cc��?�             l@������������������������       �        &             N@m       ~                    �?�qE��E�?o            �d@n       y                   �`@�q�q�?             8@o       p                   �]@      �?             0@������������������������       �                     @q       x                    r@�eP*L��?             &@r       s                    _@      �?              @������������������������       �                     �?t       w                   �m@����X�?             @u       v                   �a@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @z       {                    `P@      �?              @������������������������       �                     @|       }                    �?      �?              @������������������������       �                     �?������������������������       �                     �?       �                    �? >�֕�?[            �a@�       �                    `P@P���Q�?F            �\@�       �                    �D@ f^8���?<            �Y@�       �                   �`@����X�?             @������������������������       �                     @������������������������       �                      @�       �                   t@�q�q�?8             X@������������������������       �        1            �T@�       �                    �I@$�q-�?             *@�       �                    �H@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     $@�       �                   �j@      �?
             (@�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @�       �                    c@      �?              @������������������������       �                     @������������������������       �                     �?�       �                    �?HP�s��?             9@������������������������       �                     �?�       �                   ``@�8��8��?             8@�       �                    �M@����X�?             @�       �                   @\@�q�q�?             @������������������������       �                     �?�       �                    �F@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     1@�       �       	             �?؀�:M�?            �B@�       �                    �G@�!���?             A@������������������������       �                     &@�       �                   �j@
;&����?             7@�       �                   �`@؇���X�?             @�       �                    �M@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                 `ff�?     ��?
             0@�       �       
             �?�q�q�?             @�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @�       �                   `d@ףp=
�?             $@������������������������       �                     @�       �                 ���@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    U@���H.�?"             I@�       �                    �?ףp=
�?             4@������������������������       �                     &@�       �                 `ff�?�<ݚ�?             "@������������������������       �                     @������������������������       �                      @�       �                   pi@d��0u��?             >@������������������������       �                     @�       �                    �?
;&����?             7@������������������������       �                     @�       �                 033@ҳ�wY;�?             1@�       �                    �?և���X�?             ,@�       �                    �?؇���X�?             @�       �                 ����?r�q��?             @�       �                   0a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @r-  tr.  bh�h"h#K �r/  h%�r0  Rr1  (KK�KK�r2  hZ�Bp       �s@     0w@      p@     �]@     �l@     �Q@      (@      0@      (@                      0@     `k@      K@      1@     �C@      �?      5@      �?      @              @      �?                      1@      0@      2@       @      0@      @      �?      @              �?      �?              �?      �?              @      .@      @       @               @      @                      *@       @       @              �?       @      �?       @                      �?     @i@      .@      $@      @      "@      �?      �?      �?      �?                      �?       @              �?       @      �?                       @      h@      (@     @Q@       @      M@              &@       @      �?       @               @      �?              $@             �^@      $@      T@      "@      8@              L@      "@              @      L@      @     �G@      @     �E@      @      3@      @      3@       @      $@       @      @       @      @              @       @               @      @              @              "@                      �?      8@              @      @              @      @              "@             �E@      �?       @      �?      @              @      �?      @                      �?     �A@              ;@     �H@       @      C@              8@       @      ,@              ,@       @              9@      &@      �?      @      �?                      @      8@       @      0@      �?      &@              @      �?      @                      �?       @      @      @              @      @      @      @              @      @      �?              �?      @                      �?     �M@     �o@      C@     �k@      .@      j@              N@      .@     �b@      @      1@      @      $@              @      @      @      @      @      �?               @      @       @      �?              �?       @                      @      @              �?      @              @      �?      �?      �?                      �?       @     �`@      @     @[@      @      Y@       @      @              @       @              �?     �W@             �T@      �?      (@      �?       @               @      �?                      $@      @      "@       @       @               @       @              �?      @              @      �?               @      7@              �?       @      6@       @      @       @      �?      �?              �?      �?              �?      �?                      @              1@      7@      ,@      7@      &@      &@              (@      &@      �?      @      �?       @               @      �?                      @      &@      @       @      @       @       @       @                       @               @      "@      �?      @               @      �?       @                      �?              @      5@      =@       @      2@              &@       @      @              @       @              3@      &@      @              (@      &@      @              @      &@      @       @      @      �?      @      �?      �?      �?              �?      �?              @              �?                      @              @r3  tr4  bubhhubh)�r5  }r6  (hhh	h
hNhKhKhG        hh hNhJF<KdhG        hNhG        h@KhAKhBh"h#K �r7  h%�r8  Rr9  (KK�r:  hZ�C              �?r;  tr<  bhNh^hIC       r=  �r>  Rr?  hbKhchdKh"h#K �r@  h%�rA  RrB  (KK�rC  hI�C       rD  trE  bK�rF  RrG  }rH  (hKhnK�hoh"h#K �rI  h%�rJ  RrK  (KKυrL  hv�BH-         �                    �?bR����?�           ��@       u                   �c@2%ޑ��?           @z@       >                    �?x�����?�            x@                          �Q@��f/w�?K            �^@������������������������       �                      @       =                    �R@z�G�z�?J             ^@       <                    �?F�4�Dj�?I            �]@                        ����?��|�5��?=            �W@	                            P@�t����?             A@
                          �l@@4և���?             <@                           �?      �?             0@������������������������       �                     @                          h@8�Z$���?
             *@                          �^@�8��8��?	             (@                          `]@r�q��?             @������������������������       �                     @                          �^@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     (@                          �a@�q�q�?             @������������������������       �                     @������������������������       �                      @                        hff�?�z�G��?(             N@                           �?�<ݚ�?             "@������������������������       �                     @                          �[@���Q��?             @������������������������       �                      @������������������������       �                     @        #                    �?��[�8��?#            �I@!       "                    �?      �?             @������������������������       �                      @������������������������       �                      @$       1                    �?��k=.��?!            �G@%       0                    b@     ��?             0@&       -                    �?�q�q�?	             (@'       (                   �\@�q�q�?             "@������������������������       �                     �?)       *                   @q@      �?              @������������������������       �                     @+       ,                   0r@      �?             @������������������������       �                      @������������������������       �                      @.       /                   �m@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @2       9                    �?`Jj��?             ?@3       8                 ����? 7���B�?             ;@4       5       
             �?z�G�z�?             @������������������������       �                     �?6       7                    @K@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     6@:       ;       
             �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     8@������������������������       �                      @?       f                    �?��.���?�            pp@@       c                    `R@��ؠ���?{            `i@A       \                    �?��ֶh�?y            �h@B       [                    �M@�X�<ݺ?o            �f@C       X                    c@�[|x��?O            �_@D       E       
             �?��a��?L            @^@������������������������       �                     6@F       W                    �J@���F6��?=            �X@G       V                    �?�����H�?%            �O@H       M                    �?��a�n`�?$             O@I       J                   �a@�q�q�?             @������������������������       �                     @K       L                   �p@�q�q�?             @������������������������       �                      @������������������������       �                     �?N       O                   �U@@4և���?              L@������������������������       �                     �?P       Q                   �_@�1�`jg�?            �K@������������������������       �                    �A@R       S                    @D@R���Q�?	             4@������������������������       �                     *@T       U                   pb@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     B@Y       Z                    �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      K@]       ^                    ]@r�q��?
             2@������������������������       �                     $@_       b                    �?      �?              @`       a                   `^@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                      @d       e                    �?���Q��?             @������������������������       �                      @������������������������       �                     @g       l                   `X@�?�P�a�?'             N@h       k                    �?���Q��?             @i       j                    @K@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?m       r                    �?�C��2(�?$            �K@n       q                    �?      �?             @o       p                   �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?s       t                    �G@@9G��?             �H@������������������������       �                      @������������������������       �                    �G@v       {       
             �?��
P��?            �A@w       z                 033�?�q�q�?	             (@x       y                    �?�z�G��?             $@������������������������       �                     @������������������������       �                     @������������������������       �                      @|       }                    �?
;&����?             7@������������������������       �                     @~       �                   @b@�q�q�?
             2@       �                   m@z�G�z�?	             .@������������������������       �                     $@�       �                   0a@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                    �?�'݊U�?�            �p@�       �                   �O@�c�Α�?u            �e@�       �                   `b@ �q�q�?             8@������������������������       �                     5@�       �                    �K@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �?r�q��?g            �b@�       �                    �A@�'F����?X            �_@�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �?̌WZ�}�?V            �^@�       �       
             �?�����?H            @Z@�       �                   g@��a�n`�?             ?@������������������������       �                     @�       �                   �`@؇���X�?             <@�       �                   @[@�<ݚ�?             2@������������������������       �                     @�       �                    �G@������?             .@������������������������       �                      @�       �                   �r@8�Z$���?	             *@�       �                    �L@�8��8��?             (@������������������������       �                     "@�       �                   �_@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@�       �                   �`@xL��N�?2            �R@������������������������       �                     D@�       �                   pf@l��\��?             A@�       �                 ����?�FVQ&�?            �@@�       �                   Pb@`2U0*��?             9@������������������������       �        
             ,@�       �                   �b@�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@�       �                    a@      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                   �`@b�2�tk�?             2@�       �                   �n@և���X�?             @������������������������       �                     @������������������������       �                     @�       �                   �]@���!pc�?             &@������������������������       �                      @�       �                   �c@�����H�?             "@������������������������       �                     @�       �       	             �?�q�q�?             @�       �                    �H@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                    �?��<b���?             7@������������������������       �                     &@�       �                    @K@�q�q�?
             (@������������������������       �                     @�       �                    �?r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                    �?`�q�0ܴ?=            �W@�       �                    @L@�zvܰ?7             V@������������������������       �        0            �R@�       �                   �_@d}h���?             ,@������������������������       �                     @������������������������       �                     &@�       �                    �?r�q��?             @�       �       
             �?      �?             @�       �                     L@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @rM  trN  bh�h"h#K �rO  h%�rP  RrQ  (KK�KK�rR  hZ�B�       �q@     `y@     �P@      v@      H@     u@      :@      X@       @              8@      X@      6@      X@      6@      R@      @      >@       @      :@       @      ,@              @       @      &@      �?      &@      �?      @              @      �?      �?      �?                      �?              @      �?                      (@       @      @              @       @              2@      E@      @       @      @              @       @               @      @              &@      D@       @       @       @                       @      "@      C@      @      "@      @      @      @      @              �?      @       @      @               @       @               @       @              �?       @      �?                       @              @       @      =@      �?      :@      �?      @              �?      �?      @      �?                      @              6@      �?      @              @      �?                      8@       @              6@      n@      .@     �g@      *@      g@      $@     @e@      $@      ]@      @     �\@              6@      @      W@      @      L@      @      L@       @      @              @       @      �?       @                      �?      @      J@      �?              @      J@             �A@      @      1@              *@      @      @              @      @              �?                      B@      @       @      @                       @              K@      @      .@              $@      @      @      @      @      @                      @               @       @      @       @                      @      @     �J@       @      @       @       @               @       @                      �?      @      I@      @      @      @       @      @                       @              �?       @     �G@       @                     �G@      2@      1@      @      @      @      @      @                      @               @      &@      (@      @              @      (@      @      (@              $@      @       @      @                       @      @              k@      J@     �_@      H@      �?      7@              5@      �?       @               @      �?             @_@      9@     �Z@      4@      �?      @      �?                      @     �Z@      1@     �W@      $@      8@      @              @      8@      @      ,@      @      @              &@      @               @      &@       @      &@      �?      "@               @      �?       @                      �?              �?      $@             �Q@      @      D@              ?@      @      ?@       @      8@      �?      ,@              $@      �?              �?      $@              @      �?              �?      @                      �?      &@      @      @      @      @                      @       @      @               @       @      �?      @               @      �?      �?      �?              �?      �?              �?              2@      @      &@              @      @      @              �?      @      �?                      @     �V@      @     @U@      @     �R@              &@      @              @      &@              @      �?      @      �?      �?      �?      �?                      �?       @               @        rS  trT  bubhhubh)�rU  }rV  (hhh	h
hNhKhKhG        hh hNhJؽ�hG        hNhG        h@KhAKhBh"h#K �rW  h%�rX  RrY  (KK�rZ  hZ�C              �?r[  tr\  bhNh^hIC       r]  �r^  Rr_  hbKhchdKh"h#K �r`  h%�ra  Rrb  (KK�rc  hI�C       rd  tre  bK�rf  Rrg  }rh  (hKhnK�hoh"h#K �ri  h%�rj  Rrk  (KK��rl  hv�B�&         v                    �?z��V���?�           ��@       Y                    �?j(���?�            x@       (                    �?~�Q�$�?�             s@                           @D@V���#�?A            �W@������������������������       �                     @       '                   c@�0�~�4�?<             V@                           �?�!�,�E�?4            @R@                           �?�LQ�1	�?             7@	                          0l@���N8�?             5@
                          �a@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �        	             .@������������������������       �                      @       "                    �?H.�!���?&             I@                           �I@fP*L��?#             F@������������������������       �                     .@              	             �?>���Rp�?             =@                          �r@�J�4�?             9@                          �a@�C��2(�?             6@������������������������       �                     ,@                           X@      �?              @������������������������       �                     @                          �d@���Q��?             @������������������������       �                      @������������������������       �                     @                           �?�q�q�?             @������������������������       �                     �?                          @_@      �?              @������������������������       �                     �?������������������������       �                     �?        !                   0c@      �?             @������������������������       �                     �?������������������������       �                     @#       $                     G@�q�q�?             @������������������������       �                      @%       &                   `]@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     .@)       J                    �L@��G����?�             j@*       I                   �e@������?K            �\@+       6       
             �?��X��?J             \@,       1                    @G@؇���X�?            �A@-       0                   0b@և���X�?             @.       /                    ^@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @2       3                    �?@4և���?             <@������������������������       �                     "@4       5                    @�KM�]�?             3@������������������������       �                     1@������������������������       �                      @7       8                 ����?�kb97�?1            @S@������������������������       �                     A@9       <                    �?�ʈD��?            �E@:       ;                    _@      �?              @������������������������       �                     �?������������������������       �                     �?=       H                    �?��p\�?            �D@>       G                    j@�˹�m��?             C@?       @                   �]@      �?              @������������������������       �                      @A       B                   �\@      �?             @������������������������       �                      @C       F                   @g@      �?             @D       E                    @E@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     >@������������������������       �                     @������������������������       �                     @K       T                    c@`Ql�R�?<            �W@L       M       
             �?�|���?8             V@������������������������       �                     G@N       S                   �Z@�Ń��̧?             E@O       P                   �n@�����H�?             "@������������������������       �                     @Q       R                   �Y@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                    �@@U       X                   pc@r�q��?             @V       W                 033�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @Z       _                    �F@��}*_��?6            @T@[       \                    �?�����H�?	             2@������������������������       �                     ,@]       ^                     D@      �?             @������������������������       �                      @������������������������       �                      @`       o                   �b@�<ݚ�?-            �O@a       n                 `ff�?      �?"             H@b       i                    �?b�h�d.�?            �A@c       d                    \@�q�q�?	             (@������������������������       �                     @e       f                   @_@X�<ݚ�?             "@������������������������       �                     @g       h                   @m@�q�q�?             @������������������������       �                      @������������������������       �                     @j       k                    @M@�nkK�?             7@������������������������       �        
             *@l       m                     N@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@������������������������       �                     *@p       u                 ���@��S���?             .@q       r                   `@���!pc�?	             &@������������������������       �                     @s       t                    d@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @w       �       
             �?0�W���?�            �r@x       �                    �?(���@��?8            �W@y       z                   �a@6��f�?*            @S@������������������������       �                     >@{       |                   �e@"Ae���?            �G@������������������������       �                     "@}       �                 ���@>A�F<�?             C@~       �                    �?�MI8d�?            �B@       �                   hq@d}h���?             <@������������������������       �        
             3@�       �                    �O@�q�q�?             "@�       �                   �d@      �?              @�       �                   �r@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     "@������������������������       �                     �?�       �                    �?@�0�!��?             1@������������������������       �                     �?�       �                 033�?      �?             0@�       �                   �e@�8��8��?	             (@������������������������       �                     &@������������������������       �                     �?�       �                   �b@      �?             @������������������������       �                     @������������������������       �                     �?�       �                   Pd@� �O#�?|             j@�       �                 ����?� ��(��?y            @i@�       �                    �?�g�y��?m            @g@�       �                   `]@��Ujѡ�?>            @[@�       �                   �U@"pc�
�?             6@�       �                 ���ܿև���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �        	             .@�       �                    �M@�d���?2            �U@������������������������       �        (             R@�       �                   @\@�r����?
             .@������������������������       �                      @������������������������       �                     *@������������������������       �        /            @S@�       �                    �?     ��?             0@�       �                 ����?�q�q�?	             (@�       �                     C@�z�G��?             $@������������������������       �                      @�       �                    b@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                    �?      �?             @������������������������       �                     �?�       �                   �`@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �?؇���X�?             @������������������������       �                     �?������������������������       �                     @rm  trn  bh�h"h#K �ro  h%�rp  Rrq  (KK�KK�rr  hZ�B       pt@     �v@     �R@     `s@     �F@     0p@      ?@      P@              @      ?@     �L@      ?@      E@      4@      @      4@      �?      @      �?      @                      �?      .@                       @      &@     �C@      @     �B@              .@      @      6@      @      5@       @      4@              ,@       @      @              @       @      @       @                      @       @      �?      �?              �?      �?      �?                      �?      @      �?              �?      @              @       @       @               @       @               @       @                      .@      ,@     `h@      (@     �Y@      "@     �Y@      @      >@      @      @      �?      @      �?                      @       @               @      :@              "@       @      1@              1@       @              @     @R@              A@      @     �C@      �?      �?              �?      �?              @      C@      @     �A@      @      @               @      @      @       @              �?      @      �?      �?      �?                      �?               @              >@              @      @               @      W@      �?     �U@              G@      �?     �D@      �?       @              @      �?       @               @      �?                     �@@      �?      @      �?      �?              �?      �?                      @      >@     �I@      0@       @      ,@               @       @               @       @              ,@     �H@      @      E@      @      =@      @      @              @      @      @      @               @      @       @                      @      �?      6@              *@      �?      "@      �?                      "@              *@       @      @       @      @      @              @      @      @                      @              @     �o@     �I@      P@      >@     �N@      0@      >@              ?@      0@              "@      ?@      @      ?@      @      6@      @      3@              @      @       @      @       @       @               @       @                      @      �?              "@                      �?      @      ,@      �?               @      ,@      �?      &@              &@      �?              �?      @              @      �?             �g@      5@     `g@      .@     �f@      @     �Y@      @      2@      @      @      @      @                      @      .@             @U@       @      R@              *@       @               @      *@             @S@              @      "@      @      @      @      @       @              �?      @              @      �?               @               @       @      �?              �?       @               @      �?              �?      @      �?                      @rs  trt  bubhhubh)�ru  }rv  (hhh	h
hNhKhKhG        hh hNhJX��vhG        hNhG        h@KhAKhBh"h#K �rw  h%�rx  Rry  (KK�rz  hZ�C              �?r{  tr|  bhNh^hIC       r}  �r~  Rr  hbKhchdKh"h#K �r�  h%�r�  Rr�  (KK�r�  hI�C       r�  tr�  bK�r�  Rr�  }r�  (hKhnK�hoh"h#K �r�  h%�r�  Rr�  (KK�r�  hv�B�4         �                    �?&�b��R�?�           ��@       %                    �?�aL�C�?           �z@                          �Q@Υf���?(            �N@������������������������       �                     @                          �a@�\��N��?%            �L@                           �?�q�q�?            �C@       
                   @[@�û��|�?             7@       	                    �?      �?             @������������������������       �                     �?������������������������       �                     @                           �?�����?             3@                          �[@�r����?             .@              
             �?      �?              @������������������������       �                     �?������������������������       �                     �?                          y@$�q-�?	             *@������������������������       �                     (@������������������������       �                     �?������������������������       �                     @                          �m@      �?	             0@������������������������       �                     &@              
             �?z�G�z�?             @                          �^@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @       "                   `c@�<ݚ�?             2@       !                   �b@      �?              @                           �p@����X�?             @              
             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?#       $                   �s@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?&       �                   0b@0<o�Ɲ�?�            �v@'       (                   �U@��P��?�            Pr@������������������������       �                      @)       `                 ����?�4>�b�?�            0r@*       [                    �? ���g=�?V            @a@+       >                 ����?r�,����?8            @V@,       =                   0a@�7��?            �C@-       8                    �?�>����?             ;@.       7                   �O@���N8�?             5@/       0                    �?�C��2(�?             &@������������������������       �                     �?1       2                   `]@ףp=
�?             $@������������������������       �                     @3       4                    V@�q�q�?             @������������������������       �                     �?5       6                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@9       <                    a@r�q��?             @:       ;                    �G@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     (@?       R                   �`@�-���?             I@@       A                 033�?����"�?             =@������������������������       �                     @B       I                    �?      �?             8@C       D                   �[@և���X�?             @������������������������       �                      @E       H                    �?���Q��?             @F       G                   `Y@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?J       O       
             �?@�0�!��?
             1@K       N                    �H@      �?              @L       M                    ^@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @P       Q                    �?�<ݚ�?             "@������������������������       �                     @������������������������       �                      @S       Z                     L@�����?             5@T       Y                    �?      �?              @U       X                   �]@���Q��?             @V       W                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     *@\       ]                    �L@@�E�x�?            �H@������������������������       �                     :@^       _                   Pz@�nkK�?             7@������������������������       �                     6@������������������������       �                     �?a       |                    �?���WC�?b             c@b       y                   Ps@@P���x�?Z            �a@c       r                    �? g�yB�?Q             `@d       e                    �?��K2��?:            �W@������������������������       �                     3@f       g                   �_@�}��L�?/            �R@������������������������       �                     F@h       i       
             �?�g�y��?             ?@������������������������       �                     $@j       q       	             �?���N8�?             5@k       p                    �?�X�<ݺ?
             2@l       o                   @g@@4և���?             ,@m       n                     @      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     $@������������������������       �                     @������������������������       �                     @s       x                    @K@��?^�k�?            �A@t       u                    @؇���X�?             @������������������������       �                     @v       w                   �n@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     <@z       {                   �s@�C��2(�?	             &@������������������������       �                     �?������������������������       �                     $@}       �                 ����?$�q-�?             *@~                          �[@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     $@�       �                   d@�r*e���?/            �R@�       �                   �b@R�}e�.�?             J@�       �                 ����?؀�:M�?            �B@������������������������       �                     @�       �                    �?     ��?             @@�       �                   Pc@��
ц��?             :@�       �                    �D@�<ݚ�?             2@������������������������       �                      @�       �                   Pb@      �?             0@�       �                   �`@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �?$�q-�?	             *@������������������������       �                     @�       �       
             �?r�q��?             @������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     .@�       �                   �[@8�A�0��?             6@������������������������       �                     @�       �       	             �?�E��ӭ�?             2@�       �                   0a@8�Z$���?	             *@�       �                   �\@�8��8��?             (@�       �       
             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@������������������������       �                     �?�       �                    e@���Q��?             @������������������������       �                     �?�       �                    @M@      �?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    _@D>�Q�?�            @p@�       �                    �?�û��|�?              G@�       �                    �?��
P��?            �A@�       �                   `T@� �	��?             9@������������������������       �                     &@�       �                    �?d}h���?
             ,@������������������������       �                     @�       �                    �?�z�G��?             $@������������������������       �                     @������������������������       �                     @�       �                    ^@�z�G��?             $@�       �                   �[@�<ݚ�?             "@�       �                    `Q@���Q��?             @�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                   �^@�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?�       �                   �O@2R�T9�?�            �j@�       �                    �?؇���X�?
             ,@�       �                    �?�C��2(�?             &@������������������������       �                     @�       �                   �`@      �?              @������������������������       �                     �?������������������������       �                     @�       �                    �F@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �b@��(\���?}             i@�       �                   Pd@�IєX�?t            `g@�       �       
             �?ܴD��?D            @Y@�       �                   �b@�������?             >@�       �                 833�?���N8�?             5@�       �                    �?�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?������������������������       �                     $@�       �                     C@�q�q�?             "@�       �                   �k@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �c@r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                   �_@0z�(>��?1            �Q@������������������������       �                     C@�       �                    `@�C��2(�?            �@@������������������������       �                     �?�       �                    d@      �?             @@������������������������       �                     <@�       �                   8p@      �?             @������������������������       �                      @������������������������       �                      @�       �                    `@��f�{��?0            �U@������������������������       �                    �C@�       �                   Xt@`Ql�R�?            �G@������������������������       �                     E@�       �       
             �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                   pd@�	j*D�?	             *@������������������������       �                     @�       �                   �d@X�<ݚ�?             "@������������������������       �                     @�       �                   �l@r�q��?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KK�KK�r�  hZ�B       `r@     �x@     �S@     �u@      >@      ?@              @      >@      ;@      :@      *@      ,@      "@      �?      @      �?                      @      *@      @      *@       @      �?      �?      �?                      �?      (@      �?      (@                      �?              @      (@      @      &@              �?      @      �?       @      �?                       @               @      @      ,@      @      @       @      @       @      �?              �?       @                      @      �?              �?      "@              "@      �?             �H@     �s@      6@     �p@       @              4@     �p@      0@     �^@      .@     �R@       @     �B@       @      9@      �?      4@      �?      $@              �?      �?      "@              @      �?       @              �?      �?      �?              �?      �?                      $@      �?      @      �?       @      �?                       @              @              (@      *@     �B@      &@      2@      @              @      2@      @      @               @      @       @       @       @               @       @              �?              @      ,@      �?      @      �?      �?      �?                      �?              @       @      @              @       @               @      3@       @      @       @      @       @      �?       @                      �?               @              @              *@      �?      H@              :@      �?      6@              6@      �?              @     �b@      @      a@       @     �_@      �?     @W@              3@      �?     �R@              F@      �?      >@              $@      �?      4@      �?      1@      �?      *@      �?      @      �?                      @              $@              @              @      �?      A@      �?      @              @      �?      @              @      �?                      <@      �?      $@      �?                      $@      �?      (@      �?       @      �?                       @              $@      ;@     �G@      ,@      C@      ,@      7@              @      ,@      2@      ,@      (@      ,@      @               @      ,@       @       @      �?       @                      �?      (@      �?      @              @      �?      @              �?      �?              �?      �?                       @              @              .@      *@      "@              @      *@      @      &@       @      &@      �?      �?      �?              �?      �?              $@                      �?       @      @      �?              �?      @      �?      �?              �?      �?                       @     �j@     �F@      <@      2@      2@      1@      &@      ,@              &@      &@      @      @              @      @      @                      @      @      @      @       @      @       @      @      �?      @                      �?              �?      @                      �?      $@      �?      $@                      �?     `g@      ;@       @      (@      �?      $@              @      �?      @      �?                      @      �?       @      �?                       @      g@      .@      f@      &@     �V@      $@      7@      @      4@      �?      $@      �?      $@                      �?      $@              @      @       @      �?       @                      �?      �?      @              @      �?              Q@      @      C@              >@      @              �?      >@       @      <@               @       @               @       @             @U@      �?     �C@              G@      �?      E@              @      �?              �?      @              "@      @      @              @      @              @      @      �?      �?      �?              �?      �?              @        r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ���EhG        hNhG        h@KhAKhBh"h#K �r�  h%�r�  Rr�  (KK�r�  hZ�C              �?r�  tr�  bhNh^hIC       r�  �r�  Rr�  hbKhchdKh"h#K �r�  h%�r�  Rr�  (KK�r�  hI�C       r�  tr�  bK�r�  Rr�  }r�  (hKhnK�hoh"h#K �r�  h%�r�  Rr�  (KK݅r�  hv�BX0         �                    �K@�����?�           ��@       -                   �`@B���?�            �x@                           �?�)��?U             b@       	                    �?      �?'             Q@                          �U@(N:!���?            �A@                           �?      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     ;@
              	             �?�C��2(�?            �@@                           �E@ �Cc}�?             <@                           @B@�q�q�?             @������������������������       �                     �?������������������������       �                      @                           �?`2U0*��?             9@                           �?���N8�?	             5@                          @`@�IєX�?             1@������������������������       �                     0@������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @                          Pl@h�˹�?.             S@                            E@ ���J��?            �C@                           b@r�q��?             @������������������������       �                     @                          �`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                    �@@       ,                    �?���@��?            �B@        #       
             �?b�h�d.�?            �A@!       "                   �p@����X�?             @������������������������       �                      @������������������������       �                     @$       +                 ����?؇���X�?             <@%       &                   �m@���Q��?             $@������������������������       �                     @'       *                   @_@؇���X�?             @(       )                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �        
             2@������������������������       �                      @.       q                    �?�u4k�k�?�            �o@/       j                 ���@�q�q�?q             e@0       5                    P@�E^Y�?h            `c@1       2                    �I@d}h���?	             ,@������������������������       �                     @3       4                    �?և���X�?             @������������������������       �                     @������������������������       �                     @6       ]                   �p@��|�5��?_            �a@7       P                   �d@Vd*�=�?K            �\@8       G                   `@&����?+            @P@9       F       	             �?�z�G��?             >@:       =                    �D@��H�}�?             9@;       <                    �B@z�G�z�?             @������������������������       �                     �?������������������������       �                     @>       E                 ����?      �?             4@?       D                    d@r�q��?             2@@       A                   �b@      �?             0@������������������������       �                     &@B       C                   �\@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @H       M                    �?؇���X�?            �A@I       J                 033�? 7���B�?             ;@������������������������       �                     9@K       L                    �?      �?              @������������������������       �                     �?������������������������       �                     �?N       O                   �b@      �?              @������������������������       �                     @������������������������       �                     @Q       T                   �d@��<D�m�?             �H@R       S                    �C@      �?              @������������������������       �                     �?������������������������       �                     �?U       \                   �j@`�q�0ܴ?            �G@V       W                   e@�KM�]�?             3@������������������������       �                     �?X       [                   �\@�X�<ݺ?
             2@Y       Z                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     *@������������������������       �                     <@^       i                    �?�5��?             ;@_       h                 033�?�G��l��?             5@`       c                   `r@ҳ�wY;�?             1@a       b                   Hq@�q�q�?             @������������������������       �                      @������������������������       �                     @d       e                   0a@"pc�
�?
             &@������������������������       �                     �?f       g                    �?ףp=
�?	             $@������������������������       �                     "@������������������������       �                     �?������������������������       �                     @������������������������       �                     @k       l                    �?$�q-�?	             *@������������������������       �                     @m       p                   �j@r�q��?             @n       o                   Pb@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @r                          `c@�IєX�?5            @U@s       ~                    �?���N8�?4             U@t       u                    �?���|���?             &@������������������������       �                     �?v       y                    �?�z�G��?             $@w       x                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @z       {                   0l@؇���X�?             @������������������������       �                     @|       }                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �        .            @R@������������������������       �                     �?�       �                    �?��K��?�            0r@�       �                    �?"�W1��?�            �n@�       �                    �?�d�~V��?@            @X@�       �                 pff�?�q�q�?5             U@�       �       	             �?������?             A@�       �                    �?l��
I��?             ;@�       �                   �d@�����H�?             "@������������������������       �                      @������������������������       �                     �?�       �                    �?b�2�tk�?             2@�       �                    b@r�q��?             (@�       �                 ����?�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?������������������������       �                     �?�       �                    h@r�q��?             @������������������������       �                     @�       �                   �^@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �?j�q����?             I@�       �       	             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                 033@��0{9�?            �G@�       �                    �?      �?             <@�       �       	             �?r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                 `ff�?�C��2(�?             6@������������������������       �                     1@�       �                   �[@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     3@�       �                   �l@�θ�?             *@������������������������       �                     @�       �                    �M@և���X�?             @�       �                   �`@      �?             @������������������������       �                      @�       �                   `b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �?��(
�ɳ?Z            �b@�       �                    �L@���N8�?             5@������������������������       �                     $@�       �                   @_@�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@�       �                    @M@     8�?R             `@�       �                    �?�q��/��?             G@�       �                   @X@l��\��?             A@������������������������       �                     �?�       �                    �?�FVQ&�?            �@@�       �                   @i@�8��8��?             8@�       �       
             �?"pc�
�?             &@������������������������       �                      @�       �                   �^@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @������������������������       �        	             *@������������������������       �                     "@�       �                   P`@r�q��?             (@�       �                   �o@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �        5            �T@�       �                    @O@k��9�?            �F@�       �                    �?     ��?             @@������������������������       �                      @�       �                    V@�q�q�?             8@������������������������       �                     @�       �                     N@��Q��?             4@�       �       
             �?      �?             $@������������������������       �                     @������������������������       �                     @�       �                   �o@z�G�z�?             $@�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                   Xp@8�Z$���?             *@�       �                    �?�<ݚ�?             "@�       �                   @`@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   0m@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KK�KK�r�  hZ�B�       �s@     �w@     `m@     @d@     �E@     @Y@      A@      A@      ?@      @      @      @      @                      @      ;@              @      >@      @      9@       @      �?              �?       @              �?      8@      �?      4@      �?      0@              0@      �?                      @              @              @      "@     �P@      �?      C@      �?      @              @      �?      �?              �?      �?                     �@@       @      =@      @      =@       @      @       @                      @      @      8@      @      @      @              �?      @      �?       @      �?                       @              @              2@       @              h@     �N@      \@      L@     �[@      F@      @      &@              @      @      @              @      @              [@     �@@     @X@      1@     �I@      ,@      5@      "@      0@      "@      �?      @      �?                      @      .@      @      .@      @      .@      �?      &@              @      �?      @                      �?               @               @      @              >@      @      :@      �?      9@              �?      �?      �?                      �?      @      @      @                      @      G@      @      �?      �?              �?      �?             �F@       @      1@       @              �?      1@      �?      @      �?              �?      @              *@              <@              &@      0@      &@      $@      &@      @       @      @       @                      @      "@       @              �?      "@      �?      "@                      �?              @              @      �?      (@              @      �?      @      �?      �?              �?      �?                      @      T@      @      T@      @      @      @              �?      @      @      �?       @      �?                       @      @      �?      @               @      �?       @                      �?     @R@                      �?     @S@     �j@     �I@     `h@     �F@      J@     �A@     �H@      :@       @      3@       @       @      �?       @                      �?      &@      @      $@       @      $@      �?      $@                      �?              �?      �?      @              @      �?      �?              �?      �?              @              "@     �D@       @      �?              �?       @              @      D@      @      5@      @      �?      @                      �?       @      4@              1@       @      @       @                      @              3@      $@      @      @              @      @      �?      @               @      �?      �?      �?                      �?      @              @     �a@      �?      4@              $@      �?      $@      �?                      $@      @     �^@      @     �D@      @      ?@      �?               @      ?@       @      6@       @      "@               @       @      @              @       @                      *@              "@       @      $@       @       @       @                       @               @             �T@      :@      3@      .@      1@       @              @      1@              @      @      *@      @      @              @      @               @       @       @       @       @                       @              @      &@       @      @       @      �?      �?      �?                      �?      @      �?      @                      �?      @        r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ:9)bhG        hNhG        h@KhAKhBh"h#K �r�  h%�r�  Rr�  (KK�r�  hZ�C              �?r�  tr�  bhNh^hIC       r�  �r�  Rr�  hbKhchdKh"h#K �r�  h%�r�  Rr�  (KK�r�  hI�C       r�  tr�  bK�r�  Rr�  }r�  (hKhnK�hoh"h#K �r�  h%�r�  Rr�  (KK߅r�  hv�B�0         �                    �?�T�%y��?�           ��@       U                 ����?�H=|�P�?e           ؁@                          �O@`�J�4��?�            p@                           �I@0��_��?            �J@                           �?�㙢�c�?             7@������������������������       �                     *@                          `_@���Q��?             $@������������������������       �                     @	       
                 ����؇���X�?             @������������������������       �                     �?������������������������       �                     @                           @L@(;L]n�?             >@                           �      �?	             0@������������������������       �                     @              
             �?$�q-�?             *@������������������������       �                     @                           �?�����H�?             "@������������������������       �                     @                          �Z@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        
             ,@       @                    �?t�F�}�?�            �i@       +                    �?��8��,�?i            `c@       "                 ����?��
ц��?             :@              
             �?؇���X�?             ,@                           @K@      �?              @������������������������       �                     �?������������������������       �                     �?                           �?�8��8��?	             (@������������������������       �                      @        !                    �G@      �?             @������������������������       �                     �?������������������������       �                     @#       $                   �b@r�q��?
             (@������������������������       �                     @%       &                    �?����X�?             @������������������������       �                      @'       (                     J@���Q��?             @������������������������       �                     �?)       *                   �b@      �?             @������������������������       �                     �?������������������������       �                     @,       -                   �b@Du9iH��?T             `@������������������������       �        (            �L@.       ?                    �?      �?,             R@/       8       
             �?8^s]e�?             =@0       7                     G@���Q��?	             .@1       6                    �?�q�q�?             "@2       3                    f@      �?              @������������������������       �                     @4       5                   �\@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                     @9       >                   pf@d}h���?	             ,@:       =                   @d@�8��8��?             (@;       <                   �c@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                    �E@A       L                    �?�J��%�?            �H@B       G                     L@     ��?             @@C       F                    �?�n_Y�K�?             *@D       E                     J@      �?             $@������������������������       �                     @������������������������       �                     @������������������������       �                     @H       K                    `@�}�+r��?             3@I       J                   `Y@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        
             1@M       T                    @P@j���� �?             1@N       O                    h@����X�?             ,@������������������������       �                      @P       S                    �?r�q��?
             (@Q       R                    �B@"pc�
�?	             &@������������������������       �                      @������������������������       �                     "@������������������������       �                     �?������������������������       �                     @V       �                   �c@r�d�{�?�            �s@W       t                    �?v��؈�?�            Pq@X       e                    �?�.�+��?3            �U@Y       d                    �?և���X�?             5@Z       [                   �g@     ��?             0@������������������������       �                     @\       ]                   @_@��
ц��?	             *@������������������������       �                     @^       c                    `P@���Q��?             $@_       b                   �`@      �?              @`       a                   �q@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     @f       g                   �Q@�'�`d�?$            �P@������������������������       �                      @h       i                   P`@     ��?#             P@������������������������       �                     :@j       q                    �?�����?             C@k       l                 ����?�5��?             ;@������������������������       �                     @m       n       	             �?���N8�?	             5@������������������������       �                     .@o       p                   o@r�q��?             @������������������������       �                     @������������������������       �                     �?r       s                 `ff�?�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@u       �                    �R@�!�I�*�?v            �g@v       �                    �? .2��A�?u            �g@w       �                    �?��� ��?O             _@x       y                   �V@���!pc�?             &@������������������������       �                     �?z                           �M@z�G�z�?             $@{       |                   `c@�����H�?             "@������������������������       �                     @}       ~                   @e@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                    �? d�=��?H            @\@�       �                   �[@���N8�?C            @Z@�       �       
             �?�<ݚ�?             "@�       �                 `ff�?z�G�z�?             @������������������������       �                      @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �K@      �?             @������������������������       �                     @������������������������       �                     �?�       �                 ����?      �?;             X@�       �                    �E@�IєX�?             A@������������������������       �                     �?�       �                    �?Pa�	�?            �@@������������������������       �                     ;@�       �                   �`@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                   p@0�z��?�?#             O@������������������������       �                     D@�       �                   pp@���7�?             6@������������������������       �                     �?������������������������       �        
             5@�       �       
             �?      �?              @�       �                    �J@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                   @Y@     �?&             P@�       �                   `W@���Q��?             @������������������������       �                     @������������������������       �                      @�       �                   a@P����?$            �M@������������������������       �                    �G@�       �                 ����?�8��8��?	             (@�       �                   `a@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                    �?��%��?            �B@�       �                    �?���!pc�?             6@�       �                    a@�q�q�?             (@������������������������       �                     @������������������������       �                     @�       �                   Pj@ףp=
�?             $@�       �                 033�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    �?��S�ۿ?	             .@������������������������       �                     $@�       �                    �?z�G�z�?             @������������������������       �                     @�       �                   �q@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?x�����?N            @]@�       �                    �?(�s���?:             U@������������������������       �                     @@�       �                   Pl@4��?�?#             J@�       �                 ����?�g�y��?             ?@������������������������       �                     >@������������������������       �                     �?�       �                   @m@��s����?             5@�       �                   �l@      �?             @������������������������       �                      @�       �                    �L@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    @L@�IєX�?             1@������������������������       �                     ,@�       �                   0b@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �`@4���C�?            �@@�       �                   �a@�ՙ/�?             5@�       �                    �?      �?              @������������������������       �                      @������������������������       �                     @�       �                    �?8�Z$���?             *@�       �                     D@z�G�z�?             $@������������������������       �                     �?�       �                    �K@�����H�?             "@������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �?�8��8��?             (@������������������������       �                     $@�       �                   �l@      �?              @������������������������       �                     �?������������������������       �                     �?r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KK�KK�r�  hZ�B�       �s@     pw@     �k@     �u@      c@      Z@      @      H@      @      3@              *@      @      @      @              �?      @      �?                      @      �?      =@      �?      .@              @      �?      (@              @      �?       @              @      �?      �?      �?                      �?              ,@     �b@      L@     �`@      7@      (@      ,@       @      (@      �?      �?      �?                      �?      �?      &@               @      �?      @      �?                      @      $@       @      @              @       @       @              @       @              �?      @      �?              �?      @              ^@      "@     �L@             �O@      "@      4@      "@      "@      @      @      @       @      @              @       @      @              @       @              �?              @              &@      @      &@      �?      @      �?      @                      �?       @                       @     �E@              0@     �@@      @      :@      @       @      @      @              @      @                      @      �?      2@      �?      �?              �?      �?                      1@      $@      @      $@      @               @      $@       @      "@       @               @      "@              �?                      @     �P@     �n@     �G@     �l@      :@     �N@      (@      "@      @      "@              @      @      @      @              @      @       @      @       @       @               @       @                      @       @              @              ,@      J@       @              (@      J@              :@      (@      :@      &@      0@      @              @      0@              .@      @      �?      @                      �?      �?      $@      �?                      $@      5@      e@      3@      e@      0@      [@       @      @              �?       @       @       @      �?      @              �?      �?              �?      �?                      �?       @     @Z@      @      Y@       @      @      �?      @               @      �?       @               @      �?              �?      @              @      �?              @     @W@       @      @@      �?              �?      @@              ;@      �?      @      �?                      @      �?     �N@              D@      �?      5@      �?                      5@      @      @      �?      @      �?                      @       @              @     �N@       @      @              @       @              �?      M@             �G@      �?      &@      �?      @              @      �?                       @       @              4@      1@      @      0@      @      @              @      @              �?      "@      �?      �?      �?                      �?               @      ,@      �?      $@              @      �?      @              �?      �?              �?      �?             @W@      8@     �S@      @      @@             �G@      @      >@      �?      >@                      �?      1@      @      �?      @               @      �?      �?              �?      �?              0@      �?      ,@               @      �?              �?       @              ,@      3@      *@       @       @      @       @                      @      &@       @       @       @              �?       @      �?      @               @      �?              �?       @              @              �?      &@              $@      �?      �?              �?      �?        r�  tr�  bubhhubh)�r�  }r�  (hhh	h
hNhKhKhG        hh hNhJ�BHzhG        hNhG        h@KhAKhBh"h#K �r�  h%�r�  Rr�  (KK�r�  hZ�C              �?r�  tr�  bhNh^hIC       r�  �r�  Rr�  hbKhchdKh"h#K �r�  h%�r�  Rr�  (KK�r�  hI�C       r�  tr�  bK�r�  Rr�  }r�  (hKhnK�hoh"h#K �r�  h%�r�  Rr�  (KKǅr�  hv�B�+         �                    �?�Ba��?�           ��@       s                   �c@�i��b��?�            �w@       n       	             �?���tT��?�            �u@       S                   P`@�D��:��?�            �t@       *                    �?��%c�?j            �d@              
             �?����0�?'             K@                        033�?��S���?             .@                           �?      �?              @	                        ����?؇���X�?             @
                          �b@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?                           `P@؇���X�?             @������������������������       �                     @                           �?�q�q�?             @������������������������       �                     �?                           �?      �?              @������������������������       �                     �?������������������������       �                     �?       #                   Pa@�	j*D�?            �C@                            �?���Q��?             9@                        033�?�d�����?             3@                          �p@�n_Y�K�?             *@                          �]@���!pc�?             &@������������������������       �                     @                           �?      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                     @!       "                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?$       %                    l@؇���X�?             ,@������������������������       �                     "@&       '                    @G@���Q��?             @������������������������       �                      @(       )                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @+       N                   �a@      �?C             \@,       C                   �s@�$��y��?9            @X@-       >                    �?���1j	�?3            �U@.       9                 033@`<)�+�?.            @S@/       0                    �?������?+             R@������������������������       �                     0@1       2                    �?h�����?#             L@������������������������       �                    �G@3       4                   �]@�<ݚ�?             "@������������������������       �                     �?5       6                    �K@      �?              @������������������������       �                     @7       8                    @M@�q�q�?             @������������������������       �                     �?������������������������       �                      @:       =       
             �?z�G�z�?             @;       <                   �^@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @?       B                    Y@�<ݚ�?             "@@       A                   �\@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @D       M                    �?���|���?             &@E       J                   @_@X�<ݚ�?             "@F       G                    Z@z�G�z�?             @������������������������       �                      @H       I                     @�q�q�?             @������������������������       �                     �?������������������������       �                      @K       L                    @L@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @O       R                    �?�q�q�?
             .@P       Q                 ����?X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                     @T       g                 ����?�6,r➷?l            �d@U       V                   �?�8��8��?8             U@������������������������       �                     ?@W       Z                    �?^�!~X�?$            �J@X       Y                   �a@����X�?             ,@������������������������       �                     @������������������������       �                     $@[       \       
             �?$�q-�?            �C@������������������������       �        	             ,@]       f                   �l@H%u��?             9@^       e                   �`@     ��?             0@_       `                   `c@���!pc�?	             &@������������������������       �                     @a       b                 ����?      �?             @������������������������       �                      @c       d                   `g@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     "@h       m                    �? �)���?4            @T@i       j                   0a@�8��8��?             (@������������������������       �                     @k       l       
             �?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �        -            @Q@o       r                 `ff @�θ�?             *@p       q                   �r@�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?������������������������       �                      @t       �                    �?��+��?            �B@u       |                    �G@��}*_��?             ;@v       {       	             �?�t����?             1@w       z                    �?      �?
             0@x       y                   Xp@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     *@������������������������       �                     �?}       ~                     J@z�G�z�?             $@������������������������       �                     @       �       
             �?�q�q�?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                    �?z�G�z�?             $@�       �                 ���@�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                    �?b>:�M+�?�            0s@�       �                    �?�L���?�            0p@�       �                    @L@@H�>���?�            �k@�       �                   �d@P����?j             f@������������������������       �        D            �\@�       �                    �?Hn�.P��?&             O@������������������������       �        
             1@�       �                    �?��S�ۿ?            �F@�       �                   �b@���7�?             F@�       �                    �E@ qP��B�?            �E@������������������������       �                     7@�       �                   �e@P���Q�?             4@������������������������       �                     (@�       �                    \@      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�       �                   �p@�ʈD��?            �E@�       �                   d@؇���X�?             <@�       �                   �_@P���Q�?             4@�       �                   �o@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �        
             *@�       �                    �?      �?              @������������������������       �                     @�       �                   0g@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     .@�       �                   �O@�99lMt�?            �C@������������������������       �                     ,@������������������������       �                     9@�       �                   `b@�q�q�?             H@�       �                   �j@     ��?             @@�       �                   �`@�X�<ݺ?
             2@������������������������       �                     ,@�       �       
             �?      �?             @������������������������       �                     @������������������������       �                     �?�       �                   �^@և���X�?	             ,@�       �                   �a@���!pc�?             &@�       �                    �?      �?             @������������������������       �                      @�       �                   �[@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �?     ��?
             0@�       �       
             �?�r����?	             .@�       �                   �c@      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �?�C��2(�?             &@������������������������       �                     @�       �                    a@r�q��?             @������������������������       �                     @�       �                   @l@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?r�  tr�  bh�h"h#K �r�  h%�r�  Rr�  (KK�KK�r�  hZ�Bp       t@     �v@     �O@     �s@      F@     �r@     �D@      r@     �@@     �`@      3@     �A@      @       @      @       @      @      �?       @      �?       @                      �?      @                      �?      �?      @              @      �?       @              �?      �?      �?              �?      �?              (@      ;@      $@      .@      @      ,@      @       @      @       @              @      @      @              @      @               @                      @      @      �?      @                      �?       @      (@              "@       @      @               @       @      �?              �?       @              ,@     �X@      "@      V@      @     @T@      @     �R@       @     �Q@              0@       @      K@             �G@       @      @      �?              �?      @              @      �?       @      �?                       @      �?      @      �?       @               @      �?                       @       @      @       @      �?       @                      �?              @      @      @      @      @      �?      @               @      �?       @      �?                       @      @      �?              �?      @                       @      @      $@      @      @              @      @                      @       @     �c@      @     @S@              ?@      @      G@      @      $@      @                      $@      @      B@              ,@      @      6@      @      *@      @       @              @      @      �?       @              �?      �?      �?                      �?              @              "@      �?      T@      �?      &@              @      �?      @              @      �?                     @Q@      @      $@      �?      $@              $@      �?               @              3@      2@      1@      $@      .@       @      .@      �?       @      �?       @                      �?      *@                      �?       @       @              @       @      �?      �?      �?      �?                      �?      �?               @       @      �?       @               @      �?              �?              p@     �H@     �m@      5@     �j@      @     �e@      @     �\@             �M@      @      1@              E@      @      E@       @      E@      �?      7@              3@      �?      (@              @      �?              �?      @                      �?              �?     �C@      @      8@      @      3@      �?      @      �?      @                      �?      *@              @      @      @              �?      @      �?                      @      .@              9@      ,@              ,@      9@              4@      <@      @      9@      �?      1@              ,@      �?      @              @      �?              @       @      @       @      @      �?       @              �?      �?              �?      �?                      @      @              *@      @      *@       @      @      �?              �?      @              $@      �?      @              @      �?      @              �?      �?              �?      �?                      �?r�  tr�  bubhhubehhub.